# Copyright 2025 ICsprout Integrated Circuit Co., Ltd.
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO P65_1233_CORNER
  CLASS PAD ;
  ORIGIN 20 20 ;
  FOREIGN P65_1233_CORNER -20 -20 ;
  SIZE 130 BY 130 ;
  SYMMETRY X Y R90 ;
  SITE IOSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER MET5 ;
        RECT 99.5 103.817 107.5 110 ;
      LAYER MET4 ;
        RECT 99.5 103.817 107.5 110 ;
      LAYER MET3 ;
        RECT 99.5 103.817 107.5 110 ;
      LAYER MET2 ;
        RECT 99.5 103.817 107.5 110 ;
    END
    PORT
      LAYER MET5 ;
        RECT 103.84 99.5 110 107.5 ;
        RECT 99.5 103.817 108.75 107.504 ;
        RECT 99.5 103.817 108.742 107.531 ;
        RECT 99.5 103.817 108.696 107.577 ;
        RECT 99.5 103.817 108.65 107.623 ;
        RECT 99.5 103.817 108.604 107.669 ;
        RECT 99.5 103.817 108.558 107.715 ;
        RECT 99.5 103.817 108.512 107.761 ;
        RECT 99.5 103.817 108.466 107.807 ;
        RECT 99.5 103.817 108.42 107.853 ;
        RECT 99.5 103.817 108.374 107.899 ;
        RECT 99.5 103.817 108.328 107.945 ;
        RECT 99.5 103.817 108.282 107.991 ;
        RECT 99.5 103.817 108.236 108.037 ;
        RECT 99.5 103.817 108.19 108.083 ;
        RECT 99.5 103.817 108.144 108.129 ;
        RECT 99.5 103.817 108.098 108.175 ;
        RECT 99.5 103.817 108.052 108.221 ;
        RECT 99.5 103.817 108.006 108.267 ;
        RECT 99.5 103.817 107.96 108.313 ;
        RECT 99.5 103.817 107.914 108.359 ;
        RECT 99.5 103.817 107.868 108.405 ;
        RECT 99.5 103.817 107.822 108.451 ;
        RECT 99.5 103.817 107.776 108.497 ;
        RECT 99.5 103.817 107.73 108.543 ;
        RECT 99.5 103.817 107.684 108.589 ;
        RECT 99.5 103.817 107.638 108.635 ;
        RECT 99.5 103.817 107.592 108.681 ;
        RECT 99.5 103.817 107.546 108.727 ;
        RECT 99.546 103.771 110 107.5 ;
        RECT 103.824 99.508 107.5 110 ;
        RECT 99.592 103.725 110 107.5 ;
        RECT 103.778 99.539 107.5 110 ;
        RECT 99.638 103.679 110 107.5 ;
        RECT 103.732 99.585 107.5 110 ;
        RECT 99.684 103.633 110 107.5 ;
        RECT 103.686 99.631 107.5 110 ;
        RECT 99.73 103.587 110 107.5 ;
        RECT 103.64 99.677 107.5 110 ;
        RECT 99.776 103.541 110 107.5 ;
        RECT 103.594 99.723 107.5 110 ;
        RECT 99.822 103.495 110 107.5 ;
        RECT 103.548 99.769 107.5 110 ;
        RECT 99.868 103.449 110 107.5 ;
        RECT 103.502 99.815 107.5 110 ;
        RECT 99.914 103.403 110 107.5 ;
        RECT 103.456 99.861 107.5 110 ;
        RECT 99.96 103.357 110 107.5 ;
        RECT 103.41 99.907 107.5 110 ;
        RECT 100.006 103.311 110 107.5 ;
        RECT 103.364 99.953 107.5 110 ;
        RECT 100.052 103.265 110 107.5 ;
        RECT 103.318 99.999 107.5 110 ;
        RECT 100.098 103.219 110 107.5 ;
        RECT 103.272 100.045 107.5 110 ;
        RECT 100.144 103.173 110 107.5 ;
        RECT 103.226 100.091 107.5 110 ;
        RECT 100.19 103.127 110 107.5 ;
        RECT 103.18 100.137 107.5 110 ;
        RECT 100.236 103.081 110 107.5 ;
        RECT 103.134 100.183 107.5 110 ;
        RECT 100.282 103.035 110 107.5 ;
        RECT 103.088 100.229 107.5 110 ;
        RECT 100.328 102.989 110 107.5 ;
        RECT 103.042 100.275 107.5 110 ;
        RECT 100.374 102.943 110 107.5 ;
        RECT 102.996 100.321 107.5 110 ;
        RECT 100.42 102.897 110 107.5 ;
        RECT 102.95 100.367 107.5 110 ;
        RECT 100.466 102.851 110 107.5 ;
        RECT 102.904 100.413 107.5 110 ;
        RECT 100.512 102.805 110 107.5 ;
        RECT 102.858 100.459 107.5 110 ;
        RECT 100.558 102.759 110 107.5 ;
        RECT 102.812 100.505 107.5 110 ;
        RECT 100.604 102.713 110 107.5 ;
        RECT 102.766 100.551 107.5 110 ;
        RECT 100.65 102.667 110 107.5 ;
        RECT 102.72 100.597 107.5 110 ;
        RECT 100.696 102.621 110 107.5 ;
        RECT 102.674 100.643 107.5 110 ;
        RECT 100.742 102.575 110 107.5 ;
        RECT 102.628 100.689 107.5 110 ;
        RECT 100.788 102.529 110 107.5 ;
        RECT 102.582 100.735 107.5 110 ;
        RECT 100.834 102.483 110 107.5 ;
        RECT 102.536 100.781 107.5 110 ;
        RECT 100.88 102.437 110 107.5 ;
        RECT 102.49 100.827 107.5 110 ;
        RECT 100.926 102.391 110 107.5 ;
        RECT 102.444 100.873 107.5 110 ;
        RECT 100.972 102.345 110 107.5 ;
        RECT 102.398 100.919 107.5 110 ;
        RECT 101.018 102.299 110 107.5 ;
        RECT 102.352 100.965 107.5 110 ;
        RECT 101.064 102.253 110 107.5 ;
        RECT 102.306 101.011 107.5 110 ;
        RECT 101.11 102.207 110 107.5 ;
        RECT 102.26 101.057 107.5 110 ;
        RECT 101.156 102.161 110 107.5 ;
        RECT 102.214 101.103 107.5 110 ;
        RECT 101.202 102.115 110 107.5 ;
        RECT 102.168 101.149 107.5 110 ;
        RECT 101.248 102.069 110 107.5 ;
        RECT 102.122 101.195 107.5 110 ;
        RECT 101.294 102.023 110 107.5 ;
        RECT 102.076 101.241 107.5 110 ;
        RECT 101.34 101.977 110 107.5 ;
        RECT 102.03 101.287 107.5 110 ;
        RECT 101.386 101.931 110 107.5 ;
        RECT 101.984 101.333 107.5 110 ;
        RECT 101.432 101.885 110 107.5 ;
        RECT 101.938 101.379 107.5 110 ;
        RECT 101.478 101.839 110 107.5 ;
        RECT 101.892 101.425 107.5 110 ;
        RECT 101.524 101.793 110 107.5 ;
        RECT 101.846 101.471 107.5 110 ;
        RECT 101.57 101.747 110 107.5 ;
        RECT 101.8 101.517 107.5 110 ;
        RECT 101.616 101.701 110 107.5 ;
        RECT 101.754 101.563 107.5 110 ;
        RECT 101.662 101.655 110 107.5 ;
        RECT 101.708 101.609 107.5 110 ;
      LAYER MET4 ;
        RECT 103.84 99.5 110 107.5 ;
        RECT 99.5 103.817 108.75 107.504 ;
        RECT 99.5 103.817 108.742 107.531 ;
        RECT 99.5 103.817 108.696 107.577 ;
        RECT 99.5 103.817 108.65 107.623 ;
        RECT 99.5 103.817 108.604 107.669 ;
        RECT 99.5 103.817 108.558 107.715 ;
        RECT 99.5 103.817 108.512 107.761 ;
        RECT 99.5 103.817 108.466 107.807 ;
        RECT 99.5 103.817 108.42 107.853 ;
        RECT 99.5 103.817 108.374 107.899 ;
        RECT 99.5 103.817 108.328 107.945 ;
        RECT 99.5 103.817 108.282 107.991 ;
        RECT 99.5 103.817 108.236 108.037 ;
        RECT 99.5 103.817 108.19 108.083 ;
        RECT 99.5 103.817 108.144 108.129 ;
        RECT 99.5 103.817 108.098 108.175 ;
        RECT 99.5 103.817 108.052 108.221 ;
        RECT 99.5 103.817 108.006 108.267 ;
        RECT 99.5 103.817 107.96 108.313 ;
        RECT 99.5 103.817 107.914 108.359 ;
        RECT 99.5 103.817 107.868 108.405 ;
        RECT 99.5 103.817 107.822 108.451 ;
        RECT 99.5 103.817 107.776 108.497 ;
        RECT 99.5 103.817 107.73 108.543 ;
        RECT 99.5 103.817 107.684 108.589 ;
        RECT 99.5 103.817 107.638 108.635 ;
        RECT 99.5 103.817 107.592 108.681 ;
        RECT 99.5 103.817 107.546 108.727 ;
        RECT 99.546 103.771 110 107.5 ;
        RECT 103.824 99.508 107.5 110 ;
        RECT 99.592 103.725 110 107.5 ;
        RECT 103.778 99.539 107.5 110 ;
        RECT 99.638 103.679 110 107.5 ;
        RECT 103.732 99.585 107.5 110 ;
        RECT 99.684 103.633 110 107.5 ;
        RECT 103.686 99.631 107.5 110 ;
        RECT 99.73 103.587 110 107.5 ;
        RECT 103.64 99.677 107.5 110 ;
        RECT 99.776 103.541 110 107.5 ;
        RECT 103.594 99.723 107.5 110 ;
        RECT 99.822 103.495 110 107.5 ;
        RECT 103.548 99.769 107.5 110 ;
        RECT 99.868 103.449 110 107.5 ;
        RECT 103.502 99.815 107.5 110 ;
        RECT 99.914 103.403 110 107.5 ;
        RECT 103.456 99.861 107.5 110 ;
        RECT 99.96 103.357 110 107.5 ;
        RECT 103.41 99.907 107.5 110 ;
        RECT 100.006 103.311 110 107.5 ;
        RECT 103.364 99.953 107.5 110 ;
        RECT 100.052 103.265 110 107.5 ;
        RECT 103.318 99.999 107.5 110 ;
        RECT 100.098 103.219 110 107.5 ;
        RECT 103.272 100.045 107.5 110 ;
        RECT 100.144 103.173 110 107.5 ;
        RECT 103.226 100.091 107.5 110 ;
        RECT 100.19 103.127 110 107.5 ;
        RECT 103.18 100.137 107.5 110 ;
        RECT 100.236 103.081 110 107.5 ;
        RECT 103.134 100.183 107.5 110 ;
        RECT 100.282 103.035 110 107.5 ;
        RECT 103.088 100.229 107.5 110 ;
        RECT 100.328 102.989 110 107.5 ;
        RECT 103.042 100.275 107.5 110 ;
        RECT 100.374 102.943 110 107.5 ;
        RECT 102.996 100.321 107.5 110 ;
        RECT 100.42 102.897 110 107.5 ;
        RECT 102.95 100.367 107.5 110 ;
        RECT 100.466 102.851 110 107.5 ;
        RECT 102.904 100.413 107.5 110 ;
        RECT 100.512 102.805 110 107.5 ;
        RECT 102.858 100.459 107.5 110 ;
        RECT 100.558 102.759 110 107.5 ;
        RECT 102.812 100.505 107.5 110 ;
        RECT 100.604 102.713 110 107.5 ;
        RECT 102.766 100.551 107.5 110 ;
        RECT 100.65 102.667 110 107.5 ;
        RECT 102.72 100.597 107.5 110 ;
        RECT 100.696 102.621 110 107.5 ;
        RECT 102.674 100.643 107.5 110 ;
        RECT 100.742 102.575 110 107.5 ;
        RECT 102.628 100.689 107.5 110 ;
        RECT 100.788 102.529 110 107.5 ;
        RECT 102.582 100.735 107.5 110 ;
        RECT 100.834 102.483 110 107.5 ;
        RECT 102.536 100.781 107.5 110 ;
        RECT 100.88 102.437 110 107.5 ;
        RECT 102.49 100.827 107.5 110 ;
        RECT 100.926 102.391 110 107.5 ;
        RECT 102.444 100.873 107.5 110 ;
        RECT 100.972 102.345 110 107.5 ;
        RECT 102.398 100.919 107.5 110 ;
        RECT 101.018 102.299 110 107.5 ;
        RECT 102.352 100.965 107.5 110 ;
        RECT 101.064 102.253 110 107.5 ;
        RECT 102.306 101.011 107.5 110 ;
        RECT 101.11 102.207 110 107.5 ;
        RECT 102.26 101.057 107.5 110 ;
        RECT 101.156 102.161 110 107.5 ;
        RECT 102.214 101.103 107.5 110 ;
        RECT 101.202 102.115 110 107.5 ;
        RECT 102.168 101.149 107.5 110 ;
        RECT 101.248 102.069 110 107.5 ;
        RECT 102.122 101.195 107.5 110 ;
        RECT 101.294 102.023 110 107.5 ;
        RECT 102.076 101.241 107.5 110 ;
        RECT 101.34 101.977 110 107.5 ;
        RECT 102.03 101.287 107.5 110 ;
        RECT 101.386 101.931 110 107.5 ;
        RECT 101.984 101.333 107.5 110 ;
        RECT 101.432 101.885 110 107.5 ;
        RECT 101.938 101.379 107.5 110 ;
        RECT 101.478 101.839 110 107.5 ;
        RECT 101.892 101.425 107.5 110 ;
        RECT 101.524 101.793 110 107.5 ;
        RECT 101.846 101.471 107.5 110 ;
        RECT 101.57 101.747 110 107.5 ;
        RECT 101.8 101.517 107.5 110 ;
        RECT 101.616 101.701 110 107.5 ;
        RECT 101.754 101.563 107.5 110 ;
        RECT 101.662 101.655 110 107.5 ;
        RECT 101.708 101.609 107.5 110 ;
      LAYER MET3 ;
        RECT 103.84 99.5 110 107.5 ;
        RECT 99.5 103.817 108.75 107.504 ;
        RECT 99.5 103.817 108.742 107.531 ;
        RECT 99.5 103.817 108.696 107.577 ;
        RECT 99.5 103.817 108.65 107.623 ;
        RECT 99.5 103.817 108.604 107.669 ;
        RECT 99.5 103.817 108.558 107.715 ;
        RECT 99.5 103.817 108.512 107.761 ;
        RECT 99.5 103.817 108.466 107.807 ;
        RECT 99.5 103.817 108.42 107.853 ;
        RECT 99.5 103.817 108.374 107.899 ;
        RECT 99.5 103.817 108.328 107.945 ;
        RECT 99.5 103.817 108.282 107.991 ;
        RECT 99.5 103.817 108.236 108.037 ;
        RECT 99.5 103.817 108.19 108.083 ;
        RECT 99.5 103.817 108.144 108.129 ;
        RECT 99.5 103.817 108.098 108.175 ;
        RECT 99.5 103.817 108.052 108.221 ;
        RECT 99.5 103.817 108.006 108.267 ;
        RECT 99.5 103.817 107.96 108.313 ;
        RECT 99.5 103.817 107.914 108.359 ;
        RECT 99.5 103.817 107.868 108.405 ;
        RECT 99.5 103.817 107.822 108.451 ;
        RECT 99.5 103.817 107.776 108.497 ;
        RECT 99.5 103.817 107.73 108.543 ;
        RECT 99.5 103.817 107.684 108.589 ;
        RECT 99.5 103.817 107.638 108.635 ;
        RECT 99.5 103.817 107.592 108.681 ;
        RECT 99.5 103.817 107.546 108.727 ;
        RECT 99.546 103.771 110 107.5 ;
        RECT 103.824 99.508 107.5 110 ;
        RECT 99.592 103.725 110 107.5 ;
        RECT 103.778 99.539 107.5 110 ;
        RECT 99.638 103.679 110 107.5 ;
        RECT 103.732 99.585 107.5 110 ;
        RECT 99.684 103.633 110 107.5 ;
        RECT 103.686 99.631 107.5 110 ;
        RECT 99.73 103.587 110 107.5 ;
        RECT 103.64 99.677 107.5 110 ;
        RECT 99.776 103.541 110 107.5 ;
        RECT 103.594 99.723 107.5 110 ;
        RECT 99.822 103.495 110 107.5 ;
        RECT 103.548 99.769 107.5 110 ;
        RECT 99.868 103.449 110 107.5 ;
        RECT 103.502 99.815 107.5 110 ;
        RECT 99.914 103.403 110 107.5 ;
        RECT 103.456 99.861 107.5 110 ;
        RECT 99.96 103.357 110 107.5 ;
        RECT 103.41 99.907 107.5 110 ;
        RECT 100.006 103.311 110 107.5 ;
        RECT 103.364 99.953 107.5 110 ;
        RECT 100.052 103.265 110 107.5 ;
        RECT 103.318 99.999 107.5 110 ;
        RECT 100.098 103.219 110 107.5 ;
        RECT 103.272 100.045 107.5 110 ;
        RECT 100.144 103.173 110 107.5 ;
        RECT 103.226 100.091 107.5 110 ;
        RECT 100.19 103.127 110 107.5 ;
        RECT 103.18 100.137 107.5 110 ;
        RECT 100.236 103.081 110 107.5 ;
        RECT 103.134 100.183 107.5 110 ;
        RECT 100.282 103.035 110 107.5 ;
        RECT 103.088 100.229 107.5 110 ;
        RECT 100.328 102.989 110 107.5 ;
        RECT 103.042 100.275 107.5 110 ;
        RECT 100.374 102.943 110 107.5 ;
        RECT 102.996 100.321 107.5 110 ;
        RECT 100.42 102.897 110 107.5 ;
        RECT 102.95 100.367 107.5 110 ;
        RECT 100.466 102.851 110 107.5 ;
        RECT 102.904 100.413 107.5 110 ;
        RECT 100.512 102.805 110 107.5 ;
        RECT 102.858 100.459 107.5 110 ;
        RECT 100.558 102.759 110 107.5 ;
        RECT 102.812 100.505 107.5 110 ;
        RECT 100.604 102.713 110 107.5 ;
        RECT 102.766 100.551 107.5 110 ;
        RECT 100.65 102.667 110 107.5 ;
        RECT 102.72 100.597 107.5 110 ;
        RECT 100.696 102.621 110 107.5 ;
        RECT 102.674 100.643 107.5 110 ;
        RECT 100.742 102.575 110 107.5 ;
        RECT 102.628 100.689 107.5 110 ;
        RECT 100.788 102.529 110 107.5 ;
        RECT 102.582 100.735 107.5 110 ;
        RECT 100.834 102.483 110 107.5 ;
        RECT 102.536 100.781 107.5 110 ;
        RECT 100.88 102.437 110 107.5 ;
        RECT 102.49 100.827 107.5 110 ;
        RECT 100.926 102.391 110 107.5 ;
        RECT 102.444 100.873 107.5 110 ;
        RECT 100.972 102.345 110 107.5 ;
        RECT 102.398 100.919 107.5 110 ;
        RECT 101.018 102.299 110 107.5 ;
        RECT 102.352 100.965 107.5 110 ;
        RECT 101.064 102.253 110 107.5 ;
        RECT 102.306 101.011 107.5 110 ;
        RECT 101.11 102.207 110 107.5 ;
        RECT 102.26 101.057 107.5 110 ;
        RECT 101.156 102.161 110 107.5 ;
        RECT 102.214 101.103 107.5 110 ;
        RECT 101.202 102.115 110 107.5 ;
        RECT 102.168 101.149 107.5 110 ;
        RECT 101.248 102.069 110 107.5 ;
        RECT 102.122 101.195 107.5 110 ;
        RECT 101.294 102.023 110 107.5 ;
        RECT 102.076 101.241 107.5 110 ;
        RECT 101.34 101.977 110 107.5 ;
        RECT 102.03 101.287 107.5 110 ;
        RECT 101.386 101.931 110 107.5 ;
        RECT 101.984 101.333 107.5 110 ;
        RECT 101.432 101.885 110 107.5 ;
        RECT 101.938 101.379 107.5 110 ;
        RECT 101.478 101.839 110 107.5 ;
        RECT 101.892 101.425 107.5 110 ;
        RECT 101.524 101.793 110 107.5 ;
        RECT 101.846 101.471 107.5 110 ;
        RECT 101.57 101.747 110 107.5 ;
        RECT 101.8 101.517 107.5 110 ;
        RECT 101.616 101.701 110 107.5 ;
        RECT 101.754 101.563 107.5 110 ;
        RECT 101.662 101.655 110 107.5 ;
        RECT 101.708 101.609 107.5 110 ;
      LAYER MET2 ;
        RECT 103.84 99.5 110 107.5 ;
        RECT 99.5 103.817 108.75 107.504 ;
        RECT 99.5 103.817 108.742 107.531 ;
        RECT 99.5 103.817 108.696 107.577 ;
        RECT 99.5 103.817 108.65 107.623 ;
        RECT 99.5 103.817 108.604 107.669 ;
        RECT 99.5 103.817 108.558 107.715 ;
        RECT 99.5 103.817 108.512 107.761 ;
        RECT 99.5 103.817 108.466 107.807 ;
        RECT 99.5 103.817 108.42 107.853 ;
        RECT 99.5 103.817 108.374 107.899 ;
        RECT 99.5 103.817 108.328 107.945 ;
        RECT 99.5 103.817 108.282 107.991 ;
        RECT 99.5 103.817 108.236 108.037 ;
        RECT 99.5 103.817 108.19 108.083 ;
        RECT 99.5 103.817 108.144 108.129 ;
        RECT 99.5 103.817 108.098 108.175 ;
        RECT 99.5 103.817 108.052 108.221 ;
        RECT 99.5 103.817 108.006 108.267 ;
        RECT 99.5 103.817 107.96 108.313 ;
        RECT 99.5 103.817 107.914 108.359 ;
        RECT 99.5 103.817 107.868 108.405 ;
        RECT 99.5 103.817 107.822 108.451 ;
        RECT 99.5 103.817 107.776 108.497 ;
        RECT 99.5 103.817 107.73 108.543 ;
        RECT 99.5 103.817 107.684 108.589 ;
        RECT 99.5 103.817 107.638 108.635 ;
        RECT 99.5 103.817 107.592 108.681 ;
        RECT 99.5 103.817 107.546 108.727 ;
        RECT 99.546 103.771 110 107.5 ;
        RECT 103.824 99.508 107.5 110 ;
        RECT 99.592 103.725 110 107.5 ;
        RECT 103.778 99.539 107.5 110 ;
        RECT 99.638 103.679 110 107.5 ;
        RECT 103.732 99.585 107.5 110 ;
        RECT 99.684 103.633 110 107.5 ;
        RECT 103.686 99.631 107.5 110 ;
        RECT 99.73 103.587 110 107.5 ;
        RECT 103.64 99.677 107.5 110 ;
        RECT 99.776 103.541 110 107.5 ;
        RECT 103.594 99.723 107.5 110 ;
        RECT 99.822 103.495 110 107.5 ;
        RECT 103.548 99.769 107.5 110 ;
        RECT 99.868 103.449 110 107.5 ;
        RECT 103.502 99.815 107.5 110 ;
        RECT 99.914 103.403 110 107.5 ;
        RECT 103.456 99.861 107.5 110 ;
        RECT 99.96 103.357 110 107.5 ;
        RECT 103.41 99.907 107.5 110 ;
        RECT 100.006 103.311 110 107.5 ;
        RECT 103.364 99.953 107.5 110 ;
        RECT 100.052 103.265 110 107.5 ;
        RECT 103.318 99.999 107.5 110 ;
        RECT 100.098 103.219 110 107.5 ;
        RECT 103.272 100.045 107.5 110 ;
        RECT 100.144 103.173 110 107.5 ;
        RECT 103.226 100.091 107.5 110 ;
        RECT 100.19 103.127 110 107.5 ;
        RECT 103.18 100.137 107.5 110 ;
        RECT 100.236 103.081 110 107.5 ;
        RECT 103.134 100.183 107.5 110 ;
        RECT 100.282 103.035 110 107.5 ;
        RECT 103.088 100.229 107.5 110 ;
        RECT 100.328 102.989 110 107.5 ;
        RECT 103.042 100.275 107.5 110 ;
        RECT 100.374 102.943 110 107.5 ;
        RECT 102.996 100.321 107.5 110 ;
        RECT 100.42 102.897 110 107.5 ;
        RECT 102.95 100.367 107.5 110 ;
        RECT 100.466 102.851 110 107.5 ;
        RECT 102.904 100.413 107.5 110 ;
        RECT 100.512 102.805 110 107.5 ;
        RECT 102.858 100.459 107.5 110 ;
        RECT 100.558 102.759 110 107.5 ;
        RECT 102.812 100.505 107.5 110 ;
        RECT 100.604 102.713 110 107.5 ;
        RECT 102.766 100.551 107.5 110 ;
        RECT 100.65 102.667 110 107.5 ;
        RECT 102.72 100.597 107.5 110 ;
        RECT 100.696 102.621 110 107.5 ;
        RECT 102.674 100.643 107.5 110 ;
        RECT 100.742 102.575 110 107.5 ;
        RECT 102.628 100.689 107.5 110 ;
        RECT 100.788 102.529 110 107.5 ;
        RECT 102.582 100.735 107.5 110 ;
        RECT 100.834 102.483 110 107.5 ;
        RECT 102.536 100.781 107.5 110 ;
        RECT 100.88 102.437 110 107.5 ;
        RECT 102.49 100.827 107.5 110 ;
        RECT 100.926 102.391 110 107.5 ;
        RECT 102.444 100.873 107.5 110 ;
        RECT 100.972 102.345 110 107.5 ;
        RECT 102.398 100.919 107.5 110 ;
        RECT 101.018 102.299 110 107.5 ;
        RECT 102.352 100.965 107.5 110 ;
        RECT 101.064 102.253 110 107.5 ;
        RECT 102.306 101.011 107.5 110 ;
        RECT 101.11 102.207 110 107.5 ;
        RECT 102.26 101.057 107.5 110 ;
        RECT 101.156 102.161 110 107.5 ;
        RECT 102.214 101.103 107.5 110 ;
        RECT 101.202 102.115 110 107.5 ;
        RECT 102.168 101.149 107.5 110 ;
        RECT 101.248 102.069 110 107.5 ;
        RECT 102.122 101.195 107.5 110 ;
        RECT 101.294 102.023 110 107.5 ;
        RECT 102.076 101.241 107.5 110 ;
        RECT 101.34 101.977 110 107.5 ;
        RECT 102.03 101.287 107.5 110 ;
        RECT 101.386 101.931 110 107.5 ;
        RECT 101.984 101.333 107.5 110 ;
        RECT 101.432 101.885 110 107.5 ;
        RECT 101.938 101.379 107.5 110 ;
        RECT 101.478 101.839 110 107.5 ;
        RECT 101.892 101.425 107.5 110 ;
        RECT 101.524 101.793 110 107.5 ;
        RECT 101.846 101.471 107.5 110 ;
        RECT 101.57 101.747 110 107.5 ;
        RECT 101.8 101.517 107.5 110 ;
        RECT 101.616 101.701 110 107.5 ;
        RECT 101.754 101.563 107.5 110 ;
        RECT 101.662 101.655 110 107.5 ;
        RECT 101.708 101.609 107.5 110 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET5 ;
        RECT 79.232 61.005 79.278 69.485 ;
        RECT 70.768 69.469 79.232 69.531 ;
        RECT 77.898 62.339 110 63.5 ;
        RECT 79.186 61.051 79.232 69.531 ;
        RECT 70.722 69.515 79.186 69.577 ;
        RECT 77.944 62.293 110 63.5 ;
        RECT 79.14 61.097 79.186 69.577 ;
        RECT 70.676 69.561 79.14 69.623 ;
        RECT 77.99 62.247 110 63.5 ;
        RECT 79.094 61.143 79.14 69.623 ;
        RECT 70.63 69.607 79.094 69.669 ;
        RECT 78.036 62.201 110 63.5 ;
        RECT 79.048 61.189 79.094 69.669 ;
        RECT 70.584 69.653 79.048 69.715 ;
        RECT 78.082 62.155 110 63.5 ;
        RECT 79.002 61.235 79.048 69.715 ;
        RECT 70.538 69.699 79.002 69.761 ;
        RECT 78.128 62.109 110 63.5 ;
        RECT 78.956 61.281 79.002 69.761 ;
        RECT 70.492 69.745 78.956 69.807 ;
        RECT 78.174 62.063 110 63.5 ;
        RECT 78.91 61.327 78.956 69.807 ;
        RECT 70.446 69.791 78.91 69.853 ;
        RECT 78.22 62.017 110 63.5 ;
        RECT 78.864 61.373 78.91 69.853 ;
        RECT 70.4 69.837 78.864 69.899 ;
        RECT 78.266 61.971 110 63.5 ;
        RECT 78.818 61.419 78.864 69.899 ;
        RECT 70.354 69.883 78.818 69.945 ;
        RECT 78.312 61.925 110 63.5 ;
        RECT 78.772 61.465 78.818 69.945 ;
        RECT 70.308 69.929 78.772 69.991 ;
        RECT 78.358 61.879 110 63.5 ;
        RECT 78.726 61.511 78.772 69.991 ;
        RECT 70.262 69.975 78.726 70.037 ;
        RECT 78.404 61.833 110 63.5 ;
        RECT 78.68 61.557 78.726 70.037 ;
        RECT 70.216 70.021 78.68 70.083 ;
        RECT 78.45 61.787 110 63.5 ;
        RECT 78.634 61.603 78.68 70.083 ;
        RECT 70.17 70.067 78.634 70.129 ;
        RECT 78.496 61.741 110 63.5 ;
        RECT 78.588 61.649 78.634 70.129 ;
        RECT 70.124 70.113 78.588 70.175 ;
        RECT 78.542 61.695 110 63.5 ;
        RECT 70.078 70.159 78.542 70.221 ;
        RECT 70.032 70.205 78.496 70.267 ;
        RECT 69.986 70.251 78.45 70.313 ;
        RECT 69.94 70.297 78.404 70.359 ;
        RECT 69.894 70.343 78.358 70.405 ;
        RECT 69.848 70.389 78.312 70.451 ;
        RECT 69.802 70.435 78.266 70.497 ;
        RECT 69.756 70.481 78.22 70.543 ;
        RECT 69.71 70.527 78.174 70.589 ;
        RECT 69.664 70.573 78.128 70.635 ;
        RECT 69.618 70.619 78.082 70.681 ;
        RECT 69.572 70.665 78.036 70.727 ;
        RECT 69.526 70.711 77.99 70.773 ;
        RECT 69.48 70.757 77.944 70.819 ;
        RECT 69.434 70.803 77.898 70.865 ;
        RECT 69.388 70.849 77.852 70.911 ;
        RECT 69.342 70.895 77.806 70.957 ;
        RECT 69.296 70.941 77.76 71.003 ;
        RECT 69.25 70.987 77.714 71.049 ;
        RECT 69.204 71.033 77.668 71.095 ;
        RECT 69.158 71.079 77.622 71.141 ;
        RECT 69.112 71.125 77.576 71.187 ;
        RECT 69.066 71.171 77.53 71.233 ;
        RECT 69.02 71.217 77.484 71.279 ;
        RECT 68.974 71.263 77.438 71.325 ;
        RECT 68.928 71.309 77.392 71.371 ;
        RECT 68.882 71.355 77.346 71.417 ;
        RECT 68.836 71.401 77.3 71.463 ;
        RECT 68.79 71.447 77.254 71.509 ;
        RECT 68.744 71.493 77.208 71.555 ;
        RECT 68.698 71.539 77.162 71.601 ;
        RECT 68.652 71.585 77.116 71.647 ;
        RECT 68.606 71.631 77.07 71.693 ;
        RECT 68.56 71.677 77.024 71.739 ;
        RECT 68.514 71.723 76.978 71.785 ;
        RECT 68.468 71.769 76.932 71.831 ;
        RECT 68.422 71.815 76.886 71.877 ;
        RECT 68.376 71.861 76.84 71.923 ;
        RECT 68.33 71.907 76.794 71.969 ;
        RECT 68.284 71.953 76.748 72.015 ;
        RECT 68.238 71.999 76.702 72.061 ;
        RECT 68.192 72.045 76.656 72.107 ;
        RECT 68.146 72.091 76.61 72.153 ;
        RECT 68.1 72.137 76.564 72.199 ;
        RECT 68.054 72.183 76.518 72.245 ;
        RECT 68.008 72.229 76.472 72.291 ;
        RECT 67.962 72.275 76.426 72.337 ;
        RECT 67.916 72.321 76.38 72.383 ;
        RECT 67.87 72.367 76.334 72.429 ;
        RECT 67.824 72.413 76.288 72.475 ;
        RECT 67.778 72.459 76.242 72.521 ;
        RECT 67.732 72.505 76.196 72.567 ;
        RECT 67.686 72.551 76.15 72.613 ;
        RECT 67.64 72.597 76.104 72.659 ;
        RECT 67.594 72.643 76.058 72.705 ;
        RECT 67.548 72.689 76.012 72.751 ;
        RECT 67.502 72.735 75.966 72.797 ;
        RECT 67.456 72.781 75.92 72.843 ;
        RECT 67.41 72.827 75.874 72.889 ;
        RECT 67.364 72.873 75.828 72.935 ;
        RECT 67.318 72.919 75.782 72.981 ;
        RECT 67.272 72.965 75.736 73.027 ;
        RECT 67.226 73.011 75.69 73.073 ;
        RECT 67.18 73.057 75.644 73.119 ;
        RECT 67.134 73.103 75.598 73.165 ;
        RECT 67.088 73.149 75.552 73.211 ;
        RECT 67.042 73.195 75.506 73.257 ;
        RECT 66.996 73.241 75.46 73.303 ;
        RECT 66.95 73.287 75.414 73.349 ;
        RECT 66.904 73.333 75.368 73.395 ;
        RECT 66.858 73.379 75.322 73.441 ;
        RECT 66.812 73.425 75.276 73.487 ;
        RECT 66.766 73.471 75.23 73.533 ;
        RECT 66.72 73.517 75.184 73.579 ;
        RECT 66.674 73.563 75.138 73.625 ;
        RECT 66.628 73.609 75.092 73.671 ;
        RECT 66.582 73.655 75.046 73.717 ;
        RECT 66.536 73.701 75 73.763 ;
        RECT 66.49 73.747 74.954 73.809 ;
        RECT 66.444 73.793 74.908 73.855 ;
        RECT 66.398 73.839 74.862 73.901 ;
        RECT 66.352 73.885 74.816 73.947 ;
        RECT 66.306 73.931 74.77 73.993 ;
        RECT 66.26 73.977 74.724 74.039 ;
        RECT 66.214 74.023 74.678 74.085 ;
        RECT 66.168 74.069 74.632 74.131 ;
        RECT 66.122 74.115 74.586 74.177 ;
        RECT 66.076 74.161 74.54 74.223 ;
        RECT 66.03 74.207 74.494 74.269 ;
        RECT 65.984 74.253 74.448 74.315 ;
        RECT 65.938 74.299 74.402 74.361 ;
        RECT 65.892 74.345 74.356 74.407 ;
        RECT 65.846 74.391 74.31 74.453 ;
        RECT 65.8 74.437 74.264 74.499 ;
        RECT 65.754 74.483 74.218 74.545 ;
        RECT 65.708 74.529 74.172 74.591 ;
        RECT 65.662 74.575 74.126 74.637 ;
        RECT 65.616 74.621 74.08 74.683 ;
        RECT 65.57 74.667 74.034 74.729 ;
        RECT 65.524 74.713 73.988 74.775 ;
        RECT 65.478 74.759 73.942 74.821 ;
        RECT 65.432 74.805 73.896 74.867 ;
        RECT 65.386 74.851 73.85 74.913 ;
        RECT 65.34 74.897 73.804 74.959 ;
        RECT 65.294 74.943 73.758 75.005 ;
        RECT 65.248 74.989 73.712 75.051 ;
        RECT 65.202 75.035 73.666 75.097 ;
        RECT 65.156 75.081 73.62 75.143 ;
        RECT 65.11 75.127 73.574 75.189 ;
        RECT 65.064 75.173 73.528 75.235 ;
        RECT 65.018 75.219 73.482 75.281 ;
        RECT 64.972 75.265 73.436 75.327 ;
        RECT 64.926 75.311 73.39 75.373 ;
        RECT 64.88 75.357 73.344 75.419 ;
        RECT 64.834 75.403 73.298 75.465 ;
        RECT 64.788 75.449 73.252 75.511 ;
        RECT 64.742 75.495 73.206 75.557 ;
        RECT 64.696 75.541 73.16 75.603 ;
        RECT 64.65 75.587 73.114 75.649 ;
        RECT 64.604 75.633 73.068 75.695 ;
        RECT 64.558 75.679 73.022 75.741 ;
        RECT 64.512 75.725 72.976 75.787 ;
        RECT 64.466 75.771 72.93 75.833 ;
        RECT 64.42 75.817 72.884 75.879 ;
        RECT 64.374 75.863 72.838 75.925 ;
        RECT 64.328 75.909 72.792 75.971 ;
        RECT 64.282 75.955 72.746 76.017 ;
        RECT 64.236 76.001 72.7 76.063 ;
        RECT 64.19 76.047 72.654 76.109 ;
        RECT 64.144 76.093 72.608 76.155 ;
        RECT 64.098 76.139 72.562 76.201 ;
        RECT 64.052 76.185 72.516 76.247 ;
        RECT 64.006 76.231 72.47 76.293 ;
        RECT 63.96 76.277 72.424 76.339 ;
        RECT 63.914 76.323 72.378 76.385 ;
        RECT 63.868 76.369 72.332 76.431 ;
        RECT 63.822 76.415 72.286 76.477 ;
        RECT 63.776 76.461 72.24 76.523 ;
        RECT 63.73 76.507 72.194 76.569 ;
        RECT 63.684 76.553 72.148 76.615 ;
        RECT 63.638 76.599 72.102 76.661 ;
        RECT 63.592 76.645 72.056 76.707 ;
        RECT 63.546 76.691 72.01 76.753 ;
        RECT 63.5 76.737 71.964 76.799 ;
        RECT 63.48 76.77 71.918 76.845 ;
        RECT 63.434 76.803 71.872 76.891 ;
        RECT 63.388 76.849 71.826 76.937 ;
        RECT 63.342 76.895 71.78 76.983 ;
        RECT 63.296 76.941 71.734 77.029 ;
        RECT 63.25 76.987 71.688 77.075 ;
        RECT 63.204 77.033 71.642 77.121 ;
        RECT 63.158 77.079 71.596 77.167 ;
        RECT 63.112 77.125 71.55 77.213 ;
        RECT 63.066 77.171 71.504 77.259 ;
        RECT 63.02 77.217 71.458 77.305 ;
        RECT 62.974 77.263 71.412 77.351 ;
        RECT 62.928 77.309 71.366 77.397 ;
        RECT 62.882 77.355 71.32 77.443 ;
        RECT 62.836 77.401 71.274 77.489 ;
        RECT 62.79 77.447 71.228 77.535 ;
        RECT 62.744 77.493 71.182 77.581 ;
        RECT 62.698 77.539 71.136 77.627 ;
        RECT 62.652 77.585 71.09 77.673 ;
        RECT 62.606 77.631 71.044 77.719 ;
        RECT 62.56 77.677 70.998 77.765 ;
        RECT 62.514 77.723 70.952 77.811 ;
        RECT 62.468 77.769 70.906 77.857 ;
        RECT 62.422 77.815 70.86 77.903 ;
        RECT 62.376 77.861 70.814 77.949 ;
        RECT 62.33 77.907 70.768 77.995 ;
        RECT 62.284 77.953 70.722 78.041 ;
        RECT 62.238 77.999 70.676 78.087 ;
        RECT 62.192 78.045 70.63 78.133 ;
        RECT 62.146 78.091 70.584 78.179 ;
        RECT 62.1 78.137 70.538 78.225 ;
        RECT 62.054 78.183 70.492 78.271 ;
        RECT 62.008 78.229 70.446 78.317 ;
        RECT 61.962 78.275 70.4 78.363 ;
        RECT 61.916 78.321 70.354 78.409 ;
        RECT 61.87 78.367 70.308 78.455 ;
        RECT 61.824 78.413 70.262 78.501 ;
        RECT 61.778 78.459 70.216 78.547 ;
        RECT 61.732 78.505 70.17 78.593 ;
        RECT 61.686 78.551 70.124 78.639 ;
        RECT 61.64 78.597 70.078 78.685 ;
        RECT 61.594 78.643 70.032 78.731 ;
        RECT 61.548 78.689 69.986 78.777 ;
        RECT 61.502 78.735 69.94 78.823 ;
        RECT 61.456 78.781 69.894 78.869 ;
        RECT 61.41 78.827 69.848 78.915 ;
        RECT 61.364 78.873 69.802 78.961 ;
        RECT 61.318 78.919 69.756 79.007 ;
        RECT 61.272 78.965 69.71 79.053 ;
        RECT 61.226 79.011 69.664 79.099 ;
        RECT 61.18 79.057 69.618 79.145 ;
        RECT 61.134 79.103 69.572 79.191 ;
        RECT 61.088 79.149 69.526 79.237 ;
        RECT 61.042 79.195 69.48 79.283 ;
        RECT 60.996 79.241 69.434 79.329 ;
        RECT 60.95 79.287 69.388 79.375 ;
        RECT 60.904 79.333 69.342 79.421 ;
        RECT 60.858 79.379 69.296 79.467 ;
        RECT 60.812 79.425 69.25 79.513 ;
        RECT 60.766 79.471 69.204 79.559 ;
        RECT 60.72 79.517 69.158 79.605 ;
        RECT 60.674 79.563 69.112 79.651 ;
        RECT 60.628 79.609 69.066 79.697 ;
        RECT 60.582 79.655 69.02 79.743 ;
        RECT 60.536 79.701 68.974 79.789 ;
        RECT 60.49 79.747 68.928 79.835 ;
        RECT 60.444 79.793 68.882 79.881 ;
        RECT 60.398 79.839 68.836 79.927 ;
        RECT 60.352 79.885 68.79 79.973 ;
        RECT 60.306 79.931 68.744 80.019 ;
        RECT 60.26 79.977 68.698 80.065 ;
        RECT 60.214 80.023 68.652 80.111 ;
        RECT 60.168 80.069 68.606 80.157 ;
        RECT 60.122 80.115 68.56 80.203 ;
        RECT 60.076 80.161 68.514 80.249 ;
        RECT 60.03 80.207 68.468 80.295 ;
        RECT 59.984 80.253 68.422 80.341 ;
        RECT 59.938 80.299 68.376 80.387 ;
        RECT 59.892 80.345 68.33 80.433 ;
        RECT 59.846 80.391 68.284 80.479 ;
        RECT 59.8 80.437 68.238 80.525 ;
        RECT 59.754 80.483 68.192 80.571 ;
        RECT 59.708 80.529 68.146 80.617 ;
        RECT 59.662 80.575 68.1 80.663 ;
        RECT 59.616 80.621 68.054 80.709 ;
        RECT 59.57 80.667 68.008 80.755 ;
        RECT 59.524 80.713 67.962 80.801 ;
        RECT 59.478 80.759 67.916 80.847 ;
        RECT 59.432 80.805 67.87 80.893 ;
        RECT 59.386 80.851 67.824 80.939 ;
        RECT 59.34 80.897 67.778 80.985 ;
        RECT 59.294 80.943 67.732 81.031 ;
        RECT 59.248 80.989 67.686 81.077 ;
        RECT 59.202 81.035 67.64 81.123 ;
        RECT 59.156 81.081 67.594 81.169 ;
        RECT 59.11 81.127 67.548 81.215 ;
        RECT 59.064 81.173 67.502 81.261 ;
        RECT 59.018 81.219 67.456 81.307 ;
        RECT 58.972 81.265 67.41 81.353 ;
        RECT 58.926 81.311 67.364 81.399 ;
        RECT 58.88 81.357 67.318 81.445 ;
        RECT 58.834 81.403 67.272 81.491 ;
        RECT 58.788 81.449 67.226 81.537 ;
        RECT 58.742 81.495 67.18 81.583 ;
        RECT 58.696 81.541 67.134 81.629 ;
        RECT 58.65 81.587 67.088 81.675 ;
        RECT 58.604 81.633 67.042 81.721 ;
        RECT 58.558 81.679 66.996 81.767 ;
        RECT 58.512 81.725 66.95 81.813 ;
        RECT 58.466 81.771 66.904 81.859 ;
        RECT 58.42 81.817 66.858 81.905 ;
        RECT 58.374 81.863 66.812 81.951 ;
        RECT 58.328 81.909 66.766 81.997 ;
        RECT 58.282 81.955 66.72 82.043 ;
        RECT 58.236 82.001 66.674 82.089 ;
        RECT 58.19 82.047 66.628 82.135 ;
        RECT 58.144 82.093 66.582 82.181 ;
        RECT 58.098 82.139 66.536 82.227 ;
        RECT 58.052 82.185 66.49 82.273 ;
        RECT 58.006 82.231 66.444 82.319 ;
        RECT 57.96 82.277 66.398 82.365 ;
        RECT 57.914 82.323 66.352 82.411 ;
        RECT 57.868 82.369 66.306 82.457 ;
        RECT 57.822 82.415 66.26 82.503 ;
        RECT 57.776 82.461 66.214 82.549 ;
        RECT 57.73 82.507 66.168 82.595 ;
        RECT 57.684 82.553 66.122 82.641 ;
        RECT 57.638 82.599 66.076 82.687 ;
        RECT 57.592 82.645 66.03 82.733 ;
        RECT 57.546 82.691 65.984 82.779 ;
        RECT 57.5 82.737 65.938 82.825 ;
        RECT 57.5 82.737 65.892 82.871 ;
        RECT 57.5 82.737 65.846 82.917 ;
        RECT 57.5 82.737 65.8 82.963 ;
        RECT 57.5 82.737 65.754 83.009 ;
        RECT 57.5 82.737 65.708 83.055 ;
        RECT 57.5 82.737 65.662 83.101 ;
        RECT 57.5 82.737 65.616 83.147 ;
        RECT 57.5 82.737 65.57 83.193 ;
        RECT 57.5 82.737 65.524 83.239 ;
        RECT 57.5 82.737 65.478 83.285 ;
        RECT 57.5 82.737 65.432 83.331 ;
        RECT 57.5 82.737 65.386 83.377 ;
        RECT 57.5 82.737 65.34 83.423 ;
        RECT 57.5 82.737 65.294 83.469 ;
        RECT 57.5 82.737 65.248 83.515 ;
        RECT 57.5 82.737 65.202 83.561 ;
        RECT 57.5 82.737 65.156 83.607 ;
        RECT 57.5 82.737 65.11 83.653 ;
        RECT 57.5 82.737 65.064 83.699 ;
        RECT 57.5 82.737 65.018 83.745 ;
        RECT 57.5 82.737 64.972 83.791 ;
        RECT 57.5 82.737 64.926 83.837 ;
        RECT 57.5 82.737 64.88 83.883 ;
        RECT 57.5 82.737 64.834 83.929 ;
        RECT 57.5 82.737 64.788 83.975 ;
        RECT 57.5 82.737 64.742 84.021 ;
        RECT 57.5 82.737 64.696 84.067 ;
        RECT 57.5 82.737 64.65 84.113 ;
        RECT 57.5 82.737 64.604 84.159 ;
        RECT 57.5 82.737 64.558 84.205 ;
        RECT 57.5 82.737 64.512 84.251 ;
        RECT 57.5 82.737 64.466 84.297 ;
        RECT 57.5 82.737 64.42 84.343 ;
        RECT 57.5 82.737 64.374 84.389 ;
        RECT 57.5 82.737 64.328 84.435 ;
        RECT 57.5 82.737 64.282 84.481 ;
        RECT 57.5 82.737 64.236 84.527 ;
        RECT 57.5 82.737 64.19 84.573 ;
        RECT 57.5 82.737 64.144 84.619 ;
        RECT 57.5 82.737 64.098 84.665 ;
        RECT 57.5 82.737 64.052 84.711 ;
        RECT 57.5 82.737 64.006 84.757 ;
        RECT 57.5 82.737 63.96 84.803 ;
        RECT 57.5 82.737 63.914 84.849 ;
        RECT 57.5 82.737 63.868 84.895 ;
        RECT 57.5 82.737 63.822 84.941 ;
        RECT 57.5 82.737 63.776 84.987 ;
        RECT 57.5 82.737 63.73 85.033 ;
        RECT 57.5 82.737 63.684 85.079 ;
        RECT 57.5 82.737 63.638 85.125 ;
        RECT 57.5 82.737 63.592 85.171 ;
        RECT 57.5 82.737 63.546 85.217 ;
        RECT 57.5 82.737 63.5 110 ;
        RECT 88.365 68.5 110 77 ;
        RECT 79.852 76.99 91.885 77.012 ;
        RECT 76.366 80.476 88.365 80.522 ;
        RECT 76.412 80.43 88.411 80.497 ;
        RECT 88.362 68.501 88.365 80.522 ;
        RECT 76.458 80.384 88.457 80.451 ;
        RECT 88.316 68.526 88.362 80.546 ;
        RECT 76.32 80.522 88.316 80.592 ;
        RECT 76.504 80.338 88.503 80.405 ;
        RECT 88.27 68.572 88.316 80.592 ;
        RECT 76.274 80.568 88.27 80.638 ;
        RECT 76.55 80.292 88.549 80.359 ;
        RECT 88.224 68.618 88.27 80.638 ;
        RECT 76.228 80.614 88.224 80.684 ;
        RECT 76.596 80.246 88.595 80.313 ;
        RECT 88.178 68.664 88.224 80.684 ;
        RECT 76.182 80.66 88.178 80.73 ;
        RECT 76.642 80.2 88.641 80.267 ;
        RECT 88.132 68.71 88.178 80.73 ;
        RECT 76.136 80.706 88.132 80.776 ;
        RECT 76.688 80.154 88.687 80.221 ;
        RECT 88.086 68.756 88.132 80.776 ;
        RECT 76.09 80.752 88.086 80.822 ;
        RECT 76.734 80.108 88.733 80.175 ;
        RECT 88.04 68.802 88.086 80.822 ;
        RECT 76.044 80.798 88.04 80.868 ;
        RECT 76.78 80.062 88.779 80.129 ;
        RECT 87.994 68.848 88.04 80.868 ;
        RECT 75.998 80.844 87.994 80.914 ;
        RECT 76.826 80.016 88.825 80.083 ;
        RECT 87.948 68.894 87.994 80.914 ;
        RECT 75.952 80.89 87.948 80.96 ;
        RECT 76.872 79.97 88.871 80.037 ;
        RECT 87.902 68.94 87.948 80.96 ;
        RECT 75.906 80.936 87.902 81.006 ;
        RECT 76.918 79.924 88.917 79.991 ;
        RECT 87.856 68.986 87.902 81.006 ;
        RECT 75.86 80.982 87.856 81.052 ;
        RECT 76.964 79.883 88.963 79.945 ;
        RECT 87.81 69.032 87.856 81.052 ;
        RECT 75.814 81.028 87.81 81.098 ;
        RECT 77 79.842 89.009 79.899 ;
        RECT 87.764 69.078 87.81 81.098 ;
        RECT 75.768 81.074 87.764 81.144 ;
        RECT 77.046 79.796 89.055 79.853 ;
        RECT 87.718 69.124 87.764 81.144 ;
        RECT 75.722 81.12 87.718 81.19 ;
        RECT 77.092 79.75 89.101 79.807 ;
        RECT 87.672 69.17 87.718 81.19 ;
        RECT 75.676 81.166 87.672 81.236 ;
        RECT 77.138 79.704 89.147 79.761 ;
        RECT 87.626 69.216 87.672 81.236 ;
        RECT 75.63 81.212 87.626 81.282 ;
        RECT 77.184 79.658 89.193 79.715 ;
        RECT 87.58 69.262 87.626 81.282 ;
        RECT 75.584 81.258 87.58 81.328 ;
        RECT 77.23 79.612 89.239 79.669 ;
        RECT 87.534 69.308 87.58 81.328 ;
        RECT 75.538 81.304 87.534 81.374 ;
        RECT 77.276 79.566 89.285 79.623 ;
        RECT 87.488 69.354 87.534 81.374 ;
        RECT 75.492 81.35 87.488 81.42 ;
        RECT 77.322 79.52 89.331 79.577 ;
        RECT 87.442 69.4 87.488 81.42 ;
        RECT 75.446 81.396 87.442 81.466 ;
        RECT 77.368 79.474 89.377 79.531 ;
        RECT 87.396 69.446 87.442 81.466 ;
        RECT 75.4 81.442 87.396 81.512 ;
        RECT 77.414 79.428 89.423 79.485 ;
        RECT 87.35 69.492 87.396 81.512 ;
        RECT 75.354 81.488 87.35 81.558 ;
        RECT 77.46 79.382 89.469 79.439 ;
        RECT 87.304 69.538 87.35 81.558 ;
        RECT 75.308 81.534 87.304 81.604 ;
        RECT 77.506 79.336 89.515 79.393 ;
        RECT 87.258 69.584 87.304 81.604 ;
        RECT 75.262 81.58 87.258 81.65 ;
        RECT 77.552 79.29 89.561 79.347 ;
        RECT 87.212 69.63 87.258 81.65 ;
        RECT 75.216 81.626 87.212 81.696 ;
        RECT 77.598 79.244 89.607 79.301 ;
        RECT 87.166 69.676 87.212 81.696 ;
        RECT 75.17 81.672 87.166 81.742 ;
        RECT 77.644 79.198 89.653 79.255 ;
        RECT 87.12 69.722 87.166 81.742 ;
        RECT 75.124 81.718 87.12 81.788 ;
        RECT 77.69 79.152 89.699 79.209 ;
        RECT 87.074 69.768 87.12 81.788 ;
        RECT 75.078 81.764 87.074 81.834 ;
        RECT 77.736 79.106 89.745 79.163 ;
        RECT 87.028 69.814 87.074 81.834 ;
        RECT 75.032 81.81 87.028 81.88 ;
        RECT 77.782 79.06 89.791 79.117 ;
        RECT 86.982 69.86 87.028 81.88 ;
        RECT 74.986 81.856 86.982 81.926 ;
        RECT 77.828 79.014 89.837 79.071 ;
        RECT 86.936 69.906 86.982 81.926 ;
        RECT 74.94 81.902 86.936 81.972 ;
        RECT 77.874 78.968 89.883 79.025 ;
        RECT 86.89 69.952 86.936 81.972 ;
        RECT 74.894 81.948 86.89 82.018 ;
        RECT 77.92 78.922 89.929 78.979 ;
        RECT 86.844 69.998 86.89 82.018 ;
        RECT 74.848 81.994 86.844 82.064 ;
        RECT 77.966 78.876 89.975 78.933 ;
        RECT 86.798 70.044 86.844 82.064 ;
        RECT 74.802 82.04 86.798 82.11 ;
        RECT 78.012 78.83 90.021 78.887 ;
        RECT 86.752 70.09 86.798 82.11 ;
        RECT 74.756 82.086 86.752 82.156 ;
        RECT 78.058 78.784 90.067 78.841 ;
        RECT 86.706 70.136 86.752 82.156 ;
        RECT 74.71 82.132 86.706 82.202 ;
        RECT 78.104 78.738 90.113 78.795 ;
        RECT 86.66 70.182 86.706 82.202 ;
        RECT 74.664 82.178 86.66 82.248 ;
        RECT 78.15 78.692 90.159 78.749 ;
        RECT 86.614 70.228 86.66 82.248 ;
        RECT 74.618 82.224 86.614 82.294 ;
        RECT 78.196 78.646 90.205 78.703 ;
        RECT 86.568 70.274 86.614 82.294 ;
        RECT 74.572 82.27 86.568 82.34 ;
        RECT 78.242 78.6 90.251 78.657 ;
        RECT 86.522 70.32 86.568 82.34 ;
        RECT 74.526 82.316 86.522 82.386 ;
        RECT 78.288 78.554 90.297 78.611 ;
        RECT 86.476 70.366 86.522 82.386 ;
        RECT 74.48 82.362 86.476 82.432 ;
        RECT 78.334 78.508 90.343 78.565 ;
        RECT 86.43 70.412 86.476 82.432 ;
        RECT 74.434 82.408 86.43 82.478 ;
        RECT 78.38 78.462 90.389 78.519 ;
        RECT 86.384 70.458 86.43 82.478 ;
        RECT 74.388 82.454 86.384 82.524 ;
        RECT 78.426 78.416 90.435 78.473 ;
        RECT 86.338 70.504 86.384 82.524 ;
        RECT 74.342 82.5 86.338 82.57 ;
        RECT 78.472 78.37 90.481 78.427 ;
        RECT 86.292 70.55 86.338 82.57 ;
        RECT 74.296 82.546 86.292 82.616 ;
        RECT 78.518 78.324 90.527 78.381 ;
        RECT 86.246 70.596 86.292 82.616 ;
        RECT 74.25 82.592 86.246 82.662 ;
        RECT 78.564 78.278 90.573 78.335 ;
        RECT 86.2 70.642 86.246 82.662 ;
        RECT 74.204 82.638 86.2 82.708 ;
        RECT 78.61 78.232 90.619 78.289 ;
        RECT 86.154 70.688 86.2 82.708 ;
        RECT 74.158 82.684 86.154 82.754 ;
        RECT 78.656 78.186 90.665 78.243 ;
        RECT 86.108 70.734 86.154 82.754 ;
        RECT 74.112 82.73 86.108 82.8 ;
        RECT 78.702 78.14 90.711 78.197 ;
        RECT 86.062 70.78 86.108 82.8 ;
        RECT 74.066 82.776 86.062 82.846 ;
        RECT 78.748 78.094 90.757 78.151 ;
        RECT 86.016 70.826 86.062 82.846 ;
        RECT 74.02 82.822 86.016 82.892 ;
        RECT 78.794 78.048 90.803 78.105 ;
        RECT 85.97 70.872 86.016 82.892 ;
        RECT 73.974 82.868 85.97 82.938 ;
        RECT 78.84 78.002 90.849 78.059 ;
        RECT 85.924 70.918 85.97 82.938 ;
        RECT 73.928 82.914 85.924 82.984 ;
        RECT 78.886 77.956 90.895 78.013 ;
        RECT 85.878 70.964 85.924 82.984 ;
        RECT 73.882 82.96 85.878 83.03 ;
        RECT 78.932 77.91 90.941 77.967 ;
        RECT 85.832 71.01 85.878 83.03 ;
        RECT 73.836 83.006 85.832 83.076 ;
        RECT 78.978 77.864 90.987 77.921 ;
        RECT 85.786 71.056 85.832 83.076 ;
        RECT 73.79 83.052 85.786 83.122 ;
        RECT 79.024 77.818 91.033 77.875 ;
        RECT 85.74 71.102 85.786 83.122 ;
        RECT 73.744 83.098 85.74 83.168 ;
        RECT 79.07 77.772 91.079 77.829 ;
        RECT 85.694 71.148 85.74 83.168 ;
        RECT 73.698 83.144 85.694 83.214 ;
        RECT 79.116 77.726 91.125 77.783 ;
        RECT 85.648 71.194 85.694 83.214 ;
        RECT 73.652 83.19 85.648 83.26 ;
        RECT 79.162 77.68 91.171 77.737 ;
        RECT 85.602 71.24 85.648 83.26 ;
        RECT 73.606 83.236 85.602 83.306 ;
        RECT 79.208 77.634 91.217 77.691 ;
        RECT 85.556 71.286 85.602 83.306 ;
        RECT 73.56 83.282 85.556 83.352 ;
        RECT 79.254 77.588 91.263 77.645 ;
        RECT 85.51 71.332 85.556 83.352 ;
        RECT 73.514 83.328 85.51 83.398 ;
        RECT 79.3 77.542 91.309 77.599 ;
        RECT 85.464 71.378 85.51 83.398 ;
        RECT 73.468 83.374 85.464 83.444 ;
        RECT 79.346 77.496 91.355 77.553 ;
        RECT 85.418 71.424 85.464 83.444 ;
        RECT 73.422 83.42 85.418 83.49 ;
        RECT 79.392 77.45 91.401 77.507 ;
        RECT 85.372 71.47 85.418 83.49 ;
        RECT 73.376 83.466 85.372 83.536 ;
        RECT 79.438 77.404 91.447 77.461 ;
        RECT 85.326 71.516 85.372 83.536 ;
        RECT 73.33 83.512 85.326 83.582 ;
        RECT 79.484 77.358 91.493 77.415 ;
        RECT 85.28 71.562 85.326 83.582 ;
        RECT 73.284 83.558 85.28 83.628 ;
        RECT 79.53 77.312 91.539 77.369 ;
        RECT 85.234 71.608 85.28 83.628 ;
        RECT 73.238 83.604 85.234 83.674 ;
        RECT 79.576 77.266 91.585 77.323 ;
        RECT 85.188 71.654 85.234 83.674 ;
        RECT 73.192 83.65 85.188 83.72 ;
        RECT 79.622 77.22 91.631 77.277 ;
        RECT 85.142 71.7 85.188 83.72 ;
        RECT 73.146 83.696 85.142 83.766 ;
        RECT 79.668 77.174 91.677 77.231 ;
        RECT 85.096 71.746 85.142 83.766 ;
        RECT 73.1 83.742 85.096 83.812 ;
        RECT 79.714 77.128 91.723 77.185 ;
        RECT 85.05 71.792 85.096 83.812 ;
        RECT 73.054 83.788 85.05 83.858 ;
        RECT 79.76 77.082 91.769 77.139 ;
        RECT 85.004 71.838 85.05 83.858 ;
        RECT 73.008 83.834 85.004 83.904 ;
        RECT 79.806 77.036 91.815 77.093 ;
        RECT 84.958 71.884 85.004 83.904 ;
        RECT 72.962 83.88 84.958 83.95 ;
        RECT 79.852 76.99 91.861 77.047 ;
        RECT 84.912 71.93 84.958 83.95 ;
        RECT 72.916 83.926 84.912 83.996 ;
        RECT 79.898 76.944 110 77 ;
        RECT 84.866 71.976 84.912 83.996 ;
        RECT 72.87 83.972 84.866 84.042 ;
        RECT 79.944 76.898 110 77 ;
        RECT 84.82 72.022 84.866 84.042 ;
        RECT 72.824 84.018 84.82 84.088 ;
        RECT 79.99 76.852 110 77 ;
        RECT 84.774 72.068 84.82 84.088 ;
        RECT 72.778 84.064 84.774 84.134 ;
        RECT 80.036 76.806 110 77 ;
        RECT 84.728 72.114 84.774 84.134 ;
        RECT 72.732 84.11 84.728 84.18 ;
        RECT 80.082 76.76 110 77 ;
        RECT 84.682 72.16 84.728 84.18 ;
        RECT 72.686 84.156 84.682 84.226 ;
        RECT 80.128 76.714 110 77 ;
        RECT 84.636 72.206 84.682 84.226 ;
        RECT 72.64 84.202 84.636 84.272 ;
        RECT 80.174 76.668 110 77 ;
        RECT 84.59 72.252 84.636 84.272 ;
        RECT 72.594 84.248 84.59 84.318 ;
        RECT 80.22 76.622 110 77 ;
        RECT 84.544 72.298 84.59 84.318 ;
        RECT 72.548 84.294 84.544 84.364 ;
        RECT 80.266 76.576 110 77 ;
        RECT 84.498 72.344 84.544 84.364 ;
        RECT 72.502 84.34 84.498 84.41 ;
        RECT 80.312 76.53 110 77 ;
        RECT 84.452 72.39 84.498 84.41 ;
        RECT 72.456 84.386 84.452 84.456 ;
        RECT 80.358 76.484 110 77 ;
        RECT 84.406 72.436 84.452 84.456 ;
        RECT 72.41 84.432 84.406 84.502 ;
        RECT 80.404 76.438 110 77 ;
        RECT 84.36 72.482 84.406 84.502 ;
        RECT 72.364 84.478 84.36 84.548 ;
        RECT 80.45 76.392 110 77 ;
        RECT 84.314 72.528 84.36 84.548 ;
        RECT 72.318 84.524 84.314 84.594 ;
        RECT 80.496 76.346 110 77 ;
        RECT 84.268 72.574 84.314 84.594 ;
        RECT 72.272 84.57 84.268 84.64 ;
        RECT 80.542 76.3 110 77 ;
        RECT 84.222 72.62 84.268 84.64 ;
        RECT 72.226 84.616 84.222 84.686 ;
        RECT 80.588 76.254 110 77 ;
        RECT 84.176 72.666 84.222 84.686 ;
        RECT 72.18 84.662 84.176 84.732 ;
        RECT 80.634 76.208 110 77 ;
        RECT 84.13 72.712 84.176 84.732 ;
        RECT 72.134 84.708 84.13 84.778 ;
        RECT 80.68 76.162 110 77 ;
        RECT 84.084 72.758 84.13 84.778 ;
        RECT 72.088 84.754 84.084 84.824 ;
        RECT 80.726 76.116 110 77 ;
        RECT 84.038 72.804 84.084 84.824 ;
        RECT 72.042 84.8 84.038 84.87 ;
        RECT 80.772 76.07 110 77 ;
        RECT 83.992 72.85 84.038 84.87 ;
        RECT 71.996 84.846 83.992 84.916 ;
        RECT 80.818 76.024 110 77 ;
        RECT 83.946 72.896 83.992 84.916 ;
        RECT 71.95 84.892 83.946 84.962 ;
        RECT 80.864 75.978 110 77 ;
        RECT 83.9 72.942 83.946 84.962 ;
        RECT 71.904 84.938 83.9 85.008 ;
        RECT 80.91 75.932 110 77 ;
        RECT 83.854 72.988 83.9 85.008 ;
        RECT 71.858 84.984 83.854 85.054 ;
        RECT 80.956 75.886 110 77 ;
        RECT 83.808 73.034 83.854 85.054 ;
        RECT 71.812 85.03 83.808 85.1 ;
        RECT 81.002 75.84 110 77 ;
        RECT 83.762 73.08 83.808 85.1 ;
        RECT 71.766 85.076 83.762 85.146 ;
        RECT 81.048 75.794 110 77 ;
        RECT 83.716 73.126 83.762 85.146 ;
        RECT 71.72 85.122 83.716 85.192 ;
        RECT 81.094 75.748 110 77 ;
        RECT 83.67 73.172 83.716 85.192 ;
        RECT 71.674 85.168 83.67 85.238 ;
        RECT 81.14 75.702 110 77 ;
        RECT 83.624 73.218 83.67 85.238 ;
        RECT 71.628 85.214 83.624 85.284 ;
        RECT 81.186 75.656 110 77 ;
        RECT 83.578 73.264 83.624 85.284 ;
        RECT 71.582 85.26 83.578 85.33 ;
        RECT 81.232 75.61 110 77 ;
        RECT 83.532 73.31 83.578 85.33 ;
        RECT 71.536 85.306 83.532 85.376 ;
        RECT 81.278 75.564 110 77 ;
        RECT 83.486 73.356 83.532 85.376 ;
        RECT 71.49 85.352 83.486 85.422 ;
        RECT 81.324 75.518 110 77 ;
        RECT 83.44 73.402 83.486 85.422 ;
        RECT 71.444 85.398 83.44 85.468 ;
        RECT 81.37 75.472 110 77 ;
        RECT 83.394 73.448 83.44 85.468 ;
        RECT 71.398 85.444 83.394 85.514 ;
        RECT 81.416 75.426 110 77 ;
        RECT 83.348 73.494 83.394 85.514 ;
        RECT 71.352 85.49 83.348 85.56 ;
        RECT 81.462 75.38 110 77 ;
        RECT 83.302 73.54 83.348 85.56 ;
        RECT 71.306 85.536 83.302 85.606 ;
        RECT 81.508 75.334 110 77 ;
        RECT 83.256 73.586 83.302 85.606 ;
        RECT 71.26 85.582 83.256 85.652 ;
        RECT 81.554 75.288 110 77 ;
        RECT 83.21 73.632 83.256 85.652 ;
        RECT 71.214 85.628 83.21 85.698 ;
        RECT 81.6 75.242 110 77 ;
        RECT 83.164 73.678 83.21 85.698 ;
        RECT 71.168 85.674 83.164 85.744 ;
        RECT 81.646 75.196 110 77 ;
        RECT 83.118 73.724 83.164 85.744 ;
        RECT 71.122 85.72 83.118 85.79 ;
        RECT 81.692 75.15 110 77 ;
        RECT 83.072 73.77 83.118 85.79 ;
        RECT 71.076 85.766 83.072 85.836 ;
        RECT 81.738 75.104 110 77 ;
        RECT 83.026 73.816 83.072 85.836 ;
        RECT 71.03 85.812 83.026 85.882 ;
        RECT 81.784 75.058 110 77 ;
        RECT 82.98 73.862 83.026 85.882 ;
        RECT 70.984 85.858 82.98 85.928 ;
        RECT 81.83 75.012 110 77 ;
        RECT 82.934 73.908 82.98 85.928 ;
        RECT 70.938 85.904 82.934 85.974 ;
        RECT 81.876 74.966 110 77 ;
        RECT 82.888 73.954 82.934 85.974 ;
        RECT 70.892 85.95 82.888 86.02 ;
        RECT 81.922 74.92 110 77 ;
        RECT 82.842 74 82.888 86.02 ;
        RECT 70.846 85.996 82.842 86.066 ;
        RECT 81.968 74.874 110 77 ;
        RECT 82.796 74.046 82.842 86.066 ;
        RECT 70.8 86.042 82.796 86.112 ;
        RECT 82.014 74.828 110 77 ;
        RECT 82.75 74.092 82.796 86.112 ;
        RECT 70.754 86.088 82.75 86.158 ;
        RECT 82.06 74.782 110 77 ;
        RECT 82.704 74.138 82.75 86.158 ;
        RECT 70.708 86.134 82.704 86.204 ;
        RECT 82.106 74.736 110 77 ;
        RECT 82.658 74.184 82.704 86.204 ;
        RECT 70.662 86.18 82.658 86.25 ;
        RECT 82.152 74.69 110 77 ;
        RECT 82.612 74.23 82.658 86.25 ;
        RECT 70.616 86.226 82.612 86.296 ;
        RECT 82.198 74.644 110 77 ;
        RECT 82.566 74.276 82.612 86.296 ;
        RECT 70.57 86.272 82.566 86.342 ;
        RECT 82.244 74.598 110 77 ;
        RECT 82.52 74.322 82.566 86.342 ;
        RECT 70.524 86.318 82.52 86.388 ;
        RECT 82.29 74.552 110 77 ;
        RECT 82.474 74.368 82.52 86.388 ;
        RECT 70.478 86.364 82.474 86.434 ;
        RECT 82.336 74.506 110 77 ;
        RECT 82.428 74.414 82.474 86.434 ;
        RECT 70.432 86.41 82.428 86.48 ;
        RECT 82.382 74.46 110 77 ;
        RECT 70.386 86.456 82.382 86.526 ;
        RECT 70.34 86.502 82.336 86.572 ;
        RECT 70.294 86.548 82.29 86.618 ;
        RECT 70.248 86.594 82.244 86.664 ;
        RECT 70.202 86.64 82.198 86.71 ;
        RECT 70.156 86.686 82.152 86.756 ;
        RECT 70.11 86.732 82.106 86.802 ;
        RECT 70.064 86.778 82.06 86.848 ;
        RECT 70.018 86.824 82.014 86.894 ;
        RECT 69.972 86.87 81.968 86.94 ;
        RECT 69.926 86.916 81.922 86.986 ;
        RECT 69.88 86.962 81.876 87.032 ;
        RECT 69.834 87.008 81.83 87.078 ;
        RECT 69.788 87.054 81.784 87.124 ;
        RECT 69.742 87.1 81.738 87.17 ;
        RECT 69.696 87.146 81.692 87.216 ;
        RECT 69.65 87.192 81.646 87.262 ;
        RECT 69.604 87.238 81.6 87.308 ;
        RECT 69.558 87.284 81.554 87.354 ;
        RECT 69.512 87.33 81.508 87.4 ;
        RECT 69.466 87.376 81.462 87.446 ;
        RECT 69.42 87.422 81.416 87.492 ;
        RECT 69.374 87.468 81.37 87.538 ;
        RECT 69.328 87.514 81.324 87.584 ;
        RECT 69.282 87.56 81.278 87.63 ;
        RECT 69.236 87.606 81.232 87.676 ;
        RECT 69.19 87.652 81.186 87.722 ;
        RECT 69.144 87.698 81.14 87.768 ;
        RECT 69.098 87.744 81.094 87.814 ;
        RECT 69.052 87.79 81.048 87.86 ;
        RECT 69.006 87.836 81.002 87.906 ;
        RECT 68.96 87.882 80.956 87.952 ;
        RECT 68.914 87.928 80.91 87.998 ;
        RECT 68.868 87.974 80.864 88.044 ;
        RECT 68.822 88.02 80.818 88.09 ;
        RECT 68.776 88.066 80.772 88.136 ;
        RECT 68.73 88.112 80.726 88.182 ;
        RECT 68.684 88.158 80.68 88.228 ;
        RECT 68.638 88.204 80.634 88.274 ;
        RECT 68.592 88.25 80.588 88.32 ;
        RECT 68.546 88.296 80.542 88.366 ;
        RECT 68.5 88.342 80.496 88.412 ;
        RECT 68.5 88.342 80.45 88.458 ;
        RECT 68.5 88.342 80.404 88.504 ;
        RECT 68.5 88.342 80.358 88.55 ;
        RECT 68.5 88.342 80.312 88.596 ;
        RECT 68.5 88.342 80.266 88.642 ;
        RECT 68.5 88.342 80.22 88.688 ;
        RECT 68.5 88.342 80.174 88.734 ;
        RECT 68.5 88.342 80.128 88.78 ;
        RECT 68.5 88.342 80.082 88.826 ;
        RECT 68.5 88.342 80.036 88.872 ;
        RECT 68.5 88.342 79.99 88.918 ;
        RECT 68.5 88.342 79.944 88.964 ;
        RECT 68.5 88.342 79.898 89.01 ;
        RECT 68.5 88.342 79.852 89.056 ;
        RECT 68.5 88.342 79.806 89.102 ;
        RECT 68.5 88.342 79.76 89.148 ;
        RECT 68.5 88.342 79.714 89.194 ;
        RECT 68.5 88.342 79.668 89.24 ;
        RECT 68.5 88.342 79.622 89.286 ;
        RECT 68.5 88.342 79.576 89.332 ;
        RECT 68.5 88.342 79.53 89.378 ;
        RECT 68.5 88.342 79.484 89.424 ;
        RECT 68.5 88.342 79.438 89.47 ;
        RECT 68.5 88.342 79.392 89.516 ;
        RECT 68.5 88.342 79.346 89.562 ;
        RECT 68.5 88.342 79.3 89.608 ;
        RECT 68.5 88.342 79.254 89.654 ;
        RECT 68.5 88.342 79.208 89.7 ;
        RECT 68.5 88.342 79.162 89.746 ;
        RECT 68.5 88.342 79.116 89.792 ;
        RECT 68.5 88.342 79.07 89.838 ;
        RECT 68.5 88.342 79.024 89.884 ;
        RECT 68.5 88.342 78.978 89.93 ;
        RECT 68.5 88.342 78.932 89.976 ;
        RECT 68.5 88.342 78.886 90.022 ;
        RECT 68.5 88.342 78.84 90.068 ;
        RECT 68.5 88.342 78.794 90.114 ;
        RECT 68.5 88.342 78.748 90.16 ;
        RECT 68.5 88.342 78.702 90.206 ;
        RECT 68.5 88.342 78.656 90.252 ;
        RECT 68.5 88.342 78.61 90.298 ;
        RECT 68.5 88.342 78.564 90.344 ;
        RECT 68.5 88.342 78.518 90.39 ;
        RECT 68.5 88.342 78.472 90.436 ;
        RECT 68.5 88.342 78.426 90.482 ;
        RECT 68.5 88.342 78.38 90.528 ;
        RECT 68.5 88.342 78.334 90.574 ;
        RECT 68.5 88.342 78.288 90.62 ;
        RECT 68.5 88.342 78.242 90.666 ;
        RECT 68.5 88.342 78.196 90.712 ;
        RECT 68.5 88.342 78.15 90.758 ;
        RECT 68.5 88.342 78.104 90.804 ;
        RECT 68.5 88.342 78.058 90.85 ;
        RECT 68.5 88.342 78.012 90.896 ;
        RECT 68.5 88.342 77.966 90.942 ;
        RECT 68.5 88.342 77.92 90.988 ;
        RECT 68.5 88.342 77.874 91.034 ;
        RECT 68.5 88.342 77.828 91.08 ;
        RECT 68.5 88.342 77.782 91.126 ;
        RECT 68.5 88.342 77.736 91.172 ;
        RECT 68.5 88.342 77.69 91.218 ;
        RECT 68.5 88.342 77.644 91.264 ;
        RECT 68.5 88.342 77.598 91.31 ;
        RECT 68.5 88.342 77.552 91.356 ;
        RECT 68.5 88.342 77.506 91.402 ;
        RECT 68.5 88.342 77.46 91.448 ;
        RECT 68.5 88.342 77.414 91.494 ;
        RECT 68.5 88.342 77.368 91.54 ;
        RECT 68.5 88.342 77.322 91.586 ;
        RECT 68.5 88.342 77.276 91.632 ;
        RECT 68.5 88.342 77.23 91.678 ;
        RECT 68.5 88.342 77.184 91.724 ;
        RECT 68.5 88.342 77.138 91.77 ;
        RECT 68.5 88.342 77.092 91.816 ;
        RECT 68.5 88.342 77.046 91.862 ;
        RECT 68.5 88.342 77 110 ;
        RECT 58.714 61.528 75.642 61.611 ;
        RECT 60.002 60.24 76.955 60.298 ;
        RECT 75.596 44.646 75.642 61.611 ;
        RECT 58.668 61.574 75.596 61.657 ;
        RECT 60.048 60.194 77.001 60.252 ;
        RECT 75.55 44.692 75.596 61.657 ;
        RECT 58.622 61.62 75.55 61.703 ;
        RECT 60.094 60.148 77.047 60.206 ;
        RECT 75.504 44.738 75.55 61.703 ;
        RECT 58.576 61.666 75.504 61.749 ;
        RECT 60.14 60.102 77.093 60.16 ;
        RECT 75.458 44.784 75.504 61.749 ;
        RECT 58.53 61.712 75.458 61.795 ;
        RECT 60.186 60.056 77.139 60.114 ;
        RECT 75.412 44.83 75.458 61.795 ;
        RECT 58.484 61.758 75.412 61.841 ;
        RECT 60.232 60.01 77.185 60.068 ;
        RECT 75.366 44.876 75.412 61.841 ;
        RECT 58.438 61.804 75.366 61.887 ;
        RECT 60.278 59.964 77.231 60.022 ;
        RECT 75.32 44.922 75.366 61.887 ;
        RECT 58.392 61.85 75.32 61.933 ;
        RECT 60.324 59.918 77.277 59.976 ;
        RECT 75.274 44.968 75.32 61.933 ;
        RECT 58.346 61.896 75.274 61.979 ;
        RECT 60.37 59.872 77.323 59.93 ;
        RECT 75.228 45.014 75.274 61.979 ;
        RECT 58.3 61.942 75.228 62.025 ;
        RECT 60.416 59.826 77.369 59.884 ;
        RECT 75.182 45.06 75.228 62.025 ;
        RECT 58.254 61.988 75.182 62.071 ;
        RECT 60.462 59.78 77.415 59.838 ;
        RECT 75.136 45.106 75.182 62.071 ;
        RECT 58.208 62.034 75.136 62.117 ;
        RECT 60.508 59.734 77.461 59.792 ;
        RECT 75.09 45.152 75.136 62.117 ;
        RECT 58.162 62.08 75.09 62.163 ;
        RECT 60.554 59.688 77.507 59.746 ;
        RECT 75.044 45.198 75.09 62.163 ;
        RECT 58.116 62.126 75.044 62.209 ;
        RECT 60.6 59.642 77.553 59.7 ;
        RECT 74.998 45.244 75.044 62.209 ;
        RECT 58.07 62.172 74.998 62.255 ;
        RECT 60.646 59.596 77.599 59.654 ;
        RECT 74.952 45.29 74.998 62.255 ;
        RECT 58.024 62.218 74.952 62.301 ;
        RECT 60.692 59.55 77.645 59.608 ;
        RECT 74.906 45.336 74.952 62.301 ;
        RECT 57.978 62.264 74.906 62.347 ;
        RECT 60.738 59.504 77.691 59.562 ;
        RECT 74.86 45.382 74.906 62.347 ;
        RECT 57.932 62.31 74.86 62.393 ;
        RECT 60.784 59.458 77.737 59.516 ;
        RECT 74.814 45.428 74.86 62.393 ;
        RECT 57.886 62.356 74.814 62.439 ;
        RECT 60.83 59.412 77.783 59.47 ;
        RECT 74.768 45.474 74.814 62.439 ;
        RECT 57.84 62.402 74.768 62.485 ;
        RECT 60.876 59.366 77.829 59.424 ;
        RECT 74.722 45.52 74.768 62.485 ;
        RECT 57.794 62.448 74.722 62.531 ;
        RECT 60.922 59.32 77.875 59.378 ;
        RECT 74.676 45.566 74.722 62.531 ;
        RECT 57.748 62.494 74.676 62.577 ;
        RECT 60.968 59.274 77.921 59.332 ;
        RECT 74.63 45.612 74.676 62.577 ;
        RECT 57.702 62.54 74.63 62.623 ;
        RECT 61.014 59.228 77.967 59.286 ;
        RECT 74.584 45.658 74.63 62.623 ;
        RECT 57.656 62.586 74.584 62.669 ;
        RECT 61.06 59.182 78.013 59.24 ;
        RECT 74.538 45.704 74.584 62.669 ;
        RECT 57.61 62.632 74.538 62.715 ;
        RECT 61.106 59.136 78.059 59.194 ;
        RECT 74.492 45.75 74.538 62.715 ;
        RECT 57.564 62.678 74.492 62.761 ;
        RECT 61.152 59.09 78.105 59.148 ;
        RECT 74.446 45.796 74.492 62.761 ;
        RECT 57.518 62.724 74.446 62.807 ;
        RECT 61.198 59.044 78.151 59.102 ;
        RECT 74.4 45.842 74.446 62.807 ;
        RECT 57.472 62.77 74.4 62.853 ;
        RECT 61.244 58.998 78.197 59.056 ;
        RECT 74.354 45.888 74.4 62.853 ;
        RECT 57.426 62.816 74.354 62.899 ;
        RECT 61.29 58.952 78.243 59.01 ;
        RECT 74.308 45.934 74.354 62.899 ;
        RECT 57.38 62.862 74.308 62.945 ;
        RECT 61.336 58.906 78.289 58.964 ;
        RECT 74.262 45.98 74.308 62.945 ;
        RECT 57.334 62.908 74.262 62.991 ;
        RECT 61.382 58.86 78.335 58.918 ;
        RECT 74.216 46.026 74.262 62.991 ;
        RECT 57.288 62.954 74.216 63.037 ;
        RECT 61.428 58.814 78.381 58.872 ;
        RECT 74.17 46.072 74.216 63.037 ;
        RECT 57.242 63 74.17 63.083 ;
        RECT 61.474 58.768 78.427 58.826 ;
        RECT 74.124 46.118 74.17 63.083 ;
        RECT 57.196 63.046 74.124 63.129 ;
        RECT 61.52 58.722 78.473 58.78 ;
        RECT 74.078 46.164 74.124 63.129 ;
        RECT 57.15 63.092 74.078 63.175 ;
        RECT 61.566 58.676 78.519 58.734 ;
        RECT 74.032 46.21 74.078 63.175 ;
        RECT 57.104 63.138 74.032 63.221 ;
        RECT 61.612 58.63 78.565 58.688 ;
        RECT 73.986 46.256 74.032 63.221 ;
        RECT 57.058 63.184 73.986 63.267 ;
        RECT 61.658 58.584 78.611 58.642 ;
        RECT 73.94 46.302 73.986 63.267 ;
        RECT 57.012 63.23 73.94 63.313 ;
        RECT 61.704 58.538 78.657 58.596 ;
        RECT 73.894 46.348 73.94 63.313 ;
        RECT 56.966 63.276 73.894 63.359 ;
        RECT 61.75 58.492 78.703 58.55 ;
        RECT 73.848 46.394 73.894 63.359 ;
        RECT 56.92 63.322 73.848 63.405 ;
        RECT 61.796 58.446 78.749 58.504 ;
        RECT 73.802 46.44 73.848 63.405 ;
        RECT 56.874 63.368 73.802 63.451 ;
        RECT 61.842 58.4 78.795 58.458 ;
        RECT 73.756 46.486 73.802 63.451 ;
        RECT 56.828 63.414 73.756 63.497 ;
        RECT 61.888 58.354 78.841 58.412 ;
        RECT 73.71 46.532 73.756 63.497 ;
        RECT 56.782 63.46 73.71 63.543 ;
        RECT 61.934 58.308 78.887 58.366 ;
        RECT 73.664 46.578 73.71 63.543 ;
        RECT 56.736 63.506 73.664 63.589 ;
        RECT 61.98 58.262 78.933 58.32 ;
        RECT 73.618 46.624 73.664 63.589 ;
        RECT 56.69 63.552 73.618 63.635 ;
        RECT 62.026 58.216 78.979 58.274 ;
        RECT 73.572 46.67 73.618 63.635 ;
        RECT 56.644 63.598 73.572 63.681 ;
        RECT 62.072 58.17 79.025 58.228 ;
        RECT 73.526 46.716 73.572 63.681 ;
        RECT 56.598 63.644 73.526 63.727 ;
        RECT 62.118 58.124 79.071 58.182 ;
        RECT 73.48 46.762 73.526 63.727 ;
        RECT 56.552 63.69 73.48 63.773 ;
        RECT 62.164 58.078 79.117 58.136 ;
        RECT 73.434 46.808 73.48 63.773 ;
        RECT 56.506 63.736 73.434 63.819 ;
        RECT 62.21 58.032 79.163 58.09 ;
        RECT 73.388 46.854 73.434 63.819 ;
        RECT 56.46 63.782 73.388 63.865 ;
        RECT 62.256 57.986 79.209 58.044 ;
        RECT 73.342 46.9 73.388 63.865 ;
        RECT 56.414 63.828 73.342 63.911 ;
        RECT 62.302 57.94 79.255 57.998 ;
        RECT 73.296 46.946 73.342 63.911 ;
        RECT 56.368 63.874 73.296 63.957 ;
        RECT 62.348 57.894 79.301 57.952 ;
        RECT 73.25 46.992 73.296 63.957 ;
        RECT 56.322 63.92 73.25 64.003 ;
        RECT 62.394 57.848 79.347 57.906 ;
        RECT 73.204 47.038 73.25 64.003 ;
        RECT 56.276 63.966 73.204 64.049 ;
        RECT 62.44 57.802 79.393 57.86 ;
        RECT 73.158 47.084 73.204 64.049 ;
        RECT 56.23 64.012 73.158 64.095 ;
        RECT 62.486 57.756 79.439 57.814 ;
        RECT 73.112 47.13 73.158 64.095 ;
        RECT 56.184 64.058 73.112 64.141 ;
        RECT 62.532 57.71 79.485 57.768 ;
        RECT 73.066 47.176 73.112 64.141 ;
        RECT 56.138 64.104 73.066 64.187 ;
        RECT 62.578 57.664 79.531 57.722 ;
        RECT 73.02 47.222 73.066 64.187 ;
        RECT 56.092 64.15 73.02 64.233 ;
        RECT 62.624 57.618 79.577 57.676 ;
        RECT 72.974 47.268 73.02 64.233 ;
        RECT 56.046 64.196 72.974 64.279 ;
        RECT 62.67 57.572 79.623 57.63 ;
        RECT 72.928 47.314 72.974 64.279 ;
        RECT 56 64.242 72.928 64.325 ;
        RECT 62.716 57.526 79.669 57.584 ;
        RECT 72.882 47.36 72.928 64.325 ;
        RECT 55.96 64.285 72.882 64.371 ;
        RECT 62.762 57.48 79.715 57.538 ;
        RECT 72.836 47.406 72.882 64.371 ;
        RECT 55.914 64.328 72.836 64.417 ;
        RECT 62.808 57.434 79.761 57.492 ;
        RECT 72.79 47.452 72.836 64.417 ;
        RECT 55.868 64.374 72.79 64.463 ;
        RECT 62.854 57.388 79.807 57.446 ;
        RECT 72.744 47.498 72.79 64.463 ;
        RECT 55.822 64.42 72.744 64.509 ;
        RECT 62.9 57.342 79.853 57.4 ;
        RECT 72.698 47.544 72.744 64.509 ;
        RECT 55.776 64.466 72.698 64.555 ;
        RECT 62.946 57.296 79.899 57.354 ;
        RECT 72.652 47.59 72.698 64.555 ;
        RECT 55.73 64.512 72.652 64.601 ;
        RECT 62.992 57.25 79.945 57.308 ;
        RECT 72.606 47.636 72.652 64.601 ;
        RECT 55.684 64.558 72.606 64.647 ;
        RECT 63.038 57.204 79.991 57.262 ;
        RECT 72.56 47.682 72.606 64.647 ;
        RECT 55.638 64.604 72.56 64.693 ;
        RECT 63.084 57.158 80.037 57.216 ;
        RECT 72.514 47.728 72.56 64.693 ;
        RECT 55.592 64.65 72.514 64.739 ;
        RECT 63.13 57.112 80.083 57.17 ;
        RECT 72.468 47.774 72.514 64.739 ;
        RECT 55.546 64.696 72.468 64.785 ;
        RECT 63.176 57.066 80.129 57.124 ;
        RECT 72.422 47.82 72.468 64.785 ;
        RECT 55.5 64.742 72.422 64.831 ;
        RECT 63.222 57.02 80.175 57.078 ;
        RECT 72.376 47.866 72.422 64.831 ;
        RECT 55.454 64.788 72.376 64.877 ;
        RECT 63.268 56.974 80.221 57.032 ;
        RECT 72.33 47.912 72.376 64.877 ;
        RECT 55.408 64.834 72.33 64.923 ;
        RECT 63.314 56.928 80.267 56.986 ;
        RECT 72.284 47.958 72.33 64.923 ;
        RECT 55.362 64.88 72.284 64.969 ;
        RECT 63.36 56.882 80.313 56.94 ;
        RECT 72.238 48.004 72.284 64.969 ;
        RECT 55.316 64.926 72.238 65.015 ;
        RECT 63.406 56.836 80.359 56.894 ;
        RECT 72.192 48.05 72.238 65.015 ;
        RECT 55.27 64.972 72.192 65.061 ;
        RECT 63.452 56.79 80.405 56.848 ;
        RECT 72.146 48.096 72.192 65.061 ;
        RECT 55.224 65.018 72.146 65.107 ;
        RECT 63.498 56.744 80.451 56.802 ;
        RECT 72.1 48.142 72.146 65.107 ;
        RECT 55.178 65.064 72.1 65.153 ;
        RECT 63.544 56.698 80.497 56.756 ;
        RECT 72.054 48.188 72.1 65.153 ;
        RECT 55.132 65.11 72.054 65.199 ;
        RECT 63.59 56.652 80.543 56.71 ;
        RECT 72.008 48.234 72.054 65.199 ;
        RECT 55.086 65.156 72.008 65.245 ;
        RECT 63.636 56.606 80.589 56.664 ;
        RECT 71.962 48.28 72.008 65.245 ;
        RECT 55.04 65.202 71.962 65.291 ;
        RECT 63.682 56.56 80.635 56.618 ;
        RECT 71.916 48.326 71.962 65.291 ;
        RECT 54.994 65.248 71.916 65.337 ;
        RECT 63.728 56.514 80.681 56.572 ;
        RECT 71.87 48.372 71.916 65.337 ;
        RECT 54.948 65.294 71.87 65.383 ;
        RECT 63.774 56.468 80.727 56.526 ;
        RECT 71.824 48.418 71.87 65.383 ;
        RECT 54.902 65.34 71.824 65.429 ;
        RECT 63.82 56.422 80.773 56.48 ;
        RECT 71.778 48.464 71.824 65.429 ;
        RECT 54.856 65.386 71.778 65.475 ;
        RECT 63.866 56.376 80.819 56.434 ;
        RECT 71.732 48.51 71.778 65.475 ;
        RECT 54.81 65.432 71.732 65.521 ;
        RECT 63.912 56.33 80.865 56.388 ;
        RECT 71.686 48.556 71.732 65.521 ;
        RECT 54.764 65.478 71.686 65.567 ;
        RECT 63.958 56.284 80.911 56.342 ;
        RECT 71.64 48.602 71.686 65.567 ;
        RECT 54.718 65.524 71.64 65.613 ;
        RECT 64.004 56.238 80.957 56.296 ;
        RECT 71.594 48.648 71.64 65.613 ;
        RECT 54.672 65.57 71.594 65.659 ;
        RECT 64.05 56.192 81.003 56.25 ;
        RECT 71.548 48.694 71.594 65.659 ;
        RECT 54.626 65.616 71.548 65.705 ;
        RECT 64.096 56.146 81.049 56.204 ;
        RECT 71.502 48.74 71.548 65.705 ;
        RECT 54.58 65.662 71.502 65.751 ;
        RECT 64.142 56.1 81.095 56.158 ;
        RECT 71.456 48.786 71.502 65.751 ;
        RECT 54.534 65.708 71.456 65.797 ;
        RECT 64.188 56.054 81.141 56.112 ;
        RECT 71.41 48.832 71.456 65.797 ;
        RECT 54.488 65.754 71.41 65.843 ;
        RECT 64.234 56.008 81.187 56.066 ;
        RECT 71.364 48.878 71.41 65.843 ;
        RECT 54.442 65.8 71.364 65.889 ;
        RECT 64.28 55.962 81.23 56.022 ;
        RECT 71.318 48.924 71.364 65.889 ;
        RECT 54.396 65.846 71.318 65.935 ;
        RECT 64.326 55.916 110 56 ;
        RECT 71.272 48.97 71.318 65.935 ;
        RECT 54.35 65.892 71.272 65.981 ;
        RECT 64.372 55.87 110 56 ;
        RECT 71.226 49.016 71.272 65.981 ;
        RECT 54.304 65.938 71.226 66.027 ;
        RECT 64.418 55.824 110 56 ;
        RECT 71.18 49.062 71.226 66.027 ;
        RECT 54.258 65.984 71.18 66.073 ;
        RECT 64.464 55.778 110 56 ;
        RECT 71.134 49.108 71.18 66.073 ;
        RECT 54.212 66.03 71.134 66.119 ;
        RECT 64.51 55.732 110 56 ;
        RECT 71.088 49.154 71.134 66.119 ;
        RECT 54.166 66.076 71.088 66.165 ;
        RECT 64.556 55.686 110 56 ;
        RECT 71.042 49.2 71.088 66.165 ;
        RECT 54.12 66.122 71.042 66.211 ;
        RECT 64.602 55.64 110 56 ;
        RECT 70.996 49.246 71.042 66.211 ;
        RECT 54.074 66.168 70.996 66.257 ;
        RECT 64.648 55.594 110 56 ;
        RECT 70.95 49.292 70.996 66.257 ;
        RECT 54.028 66.214 70.95 66.303 ;
        RECT 64.694 55.548 110 56 ;
        RECT 70.904 49.338 70.95 66.303 ;
        RECT 53.982 66.26 70.904 66.349 ;
        RECT 64.74 55.502 110 56 ;
        RECT 70.858 49.384 70.904 66.349 ;
        RECT 53.936 66.306 70.858 66.395 ;
        RECT 64.786 55.456 110 56 ;
        RECT 70.812 49.43 70.858 66.395 ;
        RECT 53.89 66.352 70.812 66.441 ;
        RECT 64.832 55.41 110 56 ;
        RECT 70.766 49.476 70.812 66.441 ;
        RECT 53.844 66.398 70.766 66.487 ;
        RECT 64.878 55.364 110 56 ;
        RECT 70.72 49.522 70.766 66.487 ;
        RECT 53.798 66.444 70.72 66.533 ;
        RECT 64.924 55.318 110 56 ;
        RECT 70.674 49.568 70.72 66.533 ;
        RECT 53.752 66.49 70.674 66.579 ;
        RECT 64.97 55.272 110 56 ;
        RECT 70.628 49.614 70.674 66.579 ;
        RECT 53.706 66.536 70.628 66.625 ;
        RECT 65.016 55.226 110 56 ;
        RECT 70.582 49.66 70.628 66.625 ;
        RECT 53.66 66.582 70.582 66.671 ;
        RECT 65.062 55.18 110 56 ;
        RECT 70.536 49.706 70.582 66.671 ;
        RECT 53.614 66.628 70.536 66.717 ;
        RECT 65.108 55.134 110 56 ;
        RECT 70.49 49.752 70.536 66.717 ;
        RECT 53.568 66.674 70.49 66.763 ;
        RECT 65.154 55.088 110 56 ;
        RECT 70.444 49.798 70.49 66.763 ;
        RECT 53.522 66.72 70.444 66.809 ;
        RECT 65.2 55.042 110 56 ;
        RECT 70.398 49.844 70.444 66.809 ;
        RECT 53.476 66.766 70.398 66.855 ;
        RECT 65.246 54.996 110 56 ;
        RECT 70.352 49.89 70.398 66.855 ;
        RECT 53.43 66.812 70.352 66.901 ;
        RECT 65.292 54.95 110 56 ;
        RECT 70.306 49.936 70.352 66.901 ;
        RECT 53.384 66.858 70.306 66.947 ;
        RECT 65.338 54.904 110 56 ;
        RECT 70.26 49.982 70.306 66.947 ;
        RECT 53.338 66.904 70.26 66.993 ;
        RECT 65.384 54.858 110 56 ;
        RECT 70.214 50.028 70.26 66.993 ;
        RECT 53.292 66.95 70.214 67.039 ;
        RECT 65.43 54.812 110 56 ;
        RECT 70.168 50.074 70.214 67.039 ;
        RECT 53.246 66.996 70.168 67.085 ;
        RECT 65.476 54.766 110 56 ;
        RECT 70.122 50.12 70.168 67.085 ;
        RECT 53.2 67.042 70.122 67.131 ;
        RECT 65.522 54.72 110 56 ;
        RECT 70.076 50.166 70.122 67.131 ;
        RECT 53.154 67.088 70.076 67.177 ;
        RECT 65.568 54.674 110 56 ;
        RECT 70.03 50.212 70.076 67.177 ;
        RECT 53.108 67.134 70.03 67.223 ;
        RECT 65.614 54.628 110 56 ;
        RECT 69.984 50.258 70.03 67.223 ;
        RECT 53.062 67.18 69.984 67.269 ;
        RECT 65.66 54.582 110 56 ;
        RECT 69.938 50.304 69.984 67.269 ;
        RECT 53.016 67.226 69.938 67.315 ;
        RECT 65.706 54.536 110 56 ;
        RECT 69.892 50.35 69.938 67.315 ;
        RECT 52.97 67.272 69.892 67.361 ;
        RECT 65.752 54.49 110 56 ;
        RECT 69.846 50.396 69.892 67.361 ;
        RECT 52.924 67.318 69.846 67.407 ;
        RECT 65.798 54.444 110 56 ;
        RECT 69.8 50.442 69.846 67.407 ;
        RECT 52.878 67.364 69.8 67.453 ;
        RECT 65.844 54.398 110 56 ;
        RECT 69.754 50.488 69.8 67.453 ;
        RECT 52.832 67.41 69.754 67.499 ;
        RECT 65.89 54.352 110 56 ;
        RECT 69.708 50.534 69.754 67.499 ;
        RECT 52.786 67.456 69.708 67.545 ;
        RECT 65.936 54.306 110 56 ;
        RECT 69.662 50.58 69.708 67.545 ;
        RECT 52.74 67.502 69.662 67.591 ;
        RECT 65.982 54.26 110 56 ;
        RECT 69.616 50.626 69.662 67.591 ;
        RECT 52.694 67.548 69.616 67.637 ;
        RECT 66.028 54.214 110 56 ;
        RECT 69.57 50.672 69.616 67.637 ;
        RECT 52.648 67.594 69.57 67.683 ;
        RECT 66.074 54.168 110 56 ;
        RECT 69.524 50.718 69.57 67.683 ;
        RECT 52.602 67.64 69.524 67.729 ;
        RECT 66.12 54.122 110 56 ;
        RECT 69.478 50.764 69.524 67.729 ;
        RECT 52.556 67.686 69.478 67.775 ;
        RECT 66.166 54.076 110 56 ;
        RECT 69.432 50.81 69.478 67.775 ;
        RECT 52.51 67.732 69.432 67.821 ;
        RECT 66.212 54.03 110 56 ;
        RECT 69.386 50.856 69.432 67.821 ;
        RECT 52.464 67.778 69.386 67.867 ;
        RECT 66.258 53.984 110 56 ;
        RECT 69.34 50.902 69.386 67.867 ;
        RECT 52.418 67.824 69.34 67.913 ;
        RECT 66.304 53.938 110 56 ;
        RECT 69.294 50.948 69.34 67.913 ;
        RECT 52.372 67.87 69.294 67.959 ;
        RECT 66.35 53.892 110 56 ;
        RECT 69.248 50.994 69.294 67.959 ;
        RECT 52.326 67.916 69.248 68.005 ;
        RECT 66.396 53.846 110 56 ;
        RECT 69.202 51.04 69.248 68.005 ;
        RECT 52.28 67.962 69.202 68.051 ;
        RECT 66.442 53.8 110 56 ;
        RECT 69.156 51.086 69.202 68.051 ;
        RECT 52.234 68.008 69.156 68.097 ;
        RECT 66.488 53.754 110 56 ;
        RECT 69.11 51.132 69.156 68.097 ;
        RECT 52.188 68.054 69.11 68.143 ;
        RECT 66.534 53.708 110 56 ;
        RECT 69.064 51.178 69.11 68.143 ;
        RECT 52.142 68.1 69.064 68.189 ;
        RECT 66.58 53.662 110 56 ;
        RECT 69.018 51.224 69.064 68.189 ;
        RECT 52.096 68.146 69.018 68.235 ;
        RECT 66.626 53.616 110 56 ;
        RECT 68.972 51.27 69.018 68.235 ;
        RECT 52.05 68.192 68.972 68.281 ;
        RECT 66.672 53.57 110 56 ;
        RECT 68.926 51.316 68.972 68.281 ;
        RECT 52.004 68.238 68.926 68.327 ;
        RECT 66.718 53.524 110 56 ;
        RECT 68.88 51.362 68.926 68.327 ;
        RECT 51.958 68.284 68.88 68.373 ;
        RECT 66.764 53.478 110 56 ;
        RECT 68.834 51.408 68.88 68.373 ;
        RECT 51.912 68.33 68.834 68.419 ;
        RECT 66.81 53.432 110 56 ;
        RECT 68.788 51.454 68.834 68.419 ;
        RECT 51.866 68.376 68.788 68.465 ;
        RECT 66.856 53.386 110 56 ;
        RECT 68.742 51.5 68.788 68.465 ;
        RECT 51.82 68.422 68.742 68.511 ;
        RECT 66.902 53.34 110 56 ;
        RECT 68.696 51.546 68.742 68.511 ;
        RECT 51.774 68.468 68.696 68.557 ;
        RECT 66.948 53.294 110 56 ;
        RECT 68.65 51.592 68.696 68.557 ;
        RECT 51.728 68.514 68.65 68.603 ;
        RECT 66.994 53.248 110 56 ;
        RECT 68.604 51.638 68.65 68.603 ;
        RECT 51.682 68.56 68.604 68.649 ;
        RECT 67.04 53.202 110 56 ;
        RECT 68.558 51.684 68.604 68.649 ;
        RECT 51.636 68.606 68.558 68.695 ;
        RECT 67.086 53.156 110 56 ;
        RECT 68.512 51.73 68.558 68.695 ;
        RECT 51.59 68.652 68.512 68.741 ;
        RECT 67.132 53.11 110 56 ;
        RECT 68.466 51.776 68.512 68.741 ;
        RECT 51.544 68.698 68.466 68.787 ;
        RECT 67.178 53.064 110 56 ;
        RECT 68.42 51.822 68.466 68.787 ;
        RECT 51.498 68.744 68.42 68.833 ;
        RECT 67.224 53.018 110 56 ;
        RECT 68.374 51.868 68.42 68.833 ;
        RECT 51.452 68.79 68.374 68.879 ;
        RECT 67.27 52.972 110 56 ;
        RECT 68.328 51.914 68.374 68.879 ;
        RECT 51.406 68.836 68.328 68.925 ;
        RECT 67.316 52.926 110 56 ;
        RECT 68.282 51.96 68.328 68.925 ;
        RECT 51.36 68.882 68.282 68.971 ;
        RECT 67.362 52.88 110 56 ;
        RECT 68.236 52.006 68.282 68.971 ;
        RECT 51.314 68.928 68.236 69.017 ;
        RECT 67.408 52.834 110 56 ;
        RECT 68.19 52.052 68.236 69.017 ;
        RECT 51.268 68.974 68.19 69.063 ;
        RECT 67.454 52.788 110 56 ;
        RECT 68.144 52.098 68.19 69.063 ;
        RECT 51.222 69.02 68.144 69.109 ;
        RECT 67.5 52.742 110 56 ;
        RECT 68.098 52.144 68.144 69.109 ;
        RECT 51.176 69.066 68.098 69.155 ;
        RECT 67.546 52.696 110 56 ;
        RECT 68.052 52.19 68.098 69.155 ;
        RECT 51.13 69.112 68.052 69.201 ;
        RECT 67.592 52.65 110 56 ;
        RECT 68.006 52.236 68.052 69.201 ;
        RECT 51.084 69.158 68.006 69.247 ;
        RECT 67.638 52.604 110 56 ;
        RECT 67.96 52.282 68.006 69.247 ;
        RECT 51.038 69.204 67.96 69.293 ;
        RECT 67.684 52.558 110 56 ;
        RECT 67.914 52.328 67.96 69.293 ;
        RECT 50.992 69.25 67.914 69.339 ;
        RECT 67.73 52.512 110 56 ;
        RECT 67.868 52.374 67.914 69.339 ;
        RECT 50.946 69.296 67.868 69.385 ;
        RECT 67.776 52.466 110 56 ;
        RECT 67.822 52.42 67.868 69.385 ;
        RECT 50.9 69.342 67.822 69.431 ;
        RECT 50.854 69.388 67.776 69.477 ;
        RECT 50.808 69.434 67.73 69.523 ;
        RECT 50.762 69.48 67.684 69.569 ;
        RECT 50.716 69.526 67.638 69.615 ;
        RECT 50.67 69.572 67.592 69.661 ;
        RECT 50.624 69.618 67.546 69.707 ;
        RECT 50.578 69.664 67.5 69.753 ;
        RECT 50.532 69.71 67.454 69.799 ;
        RECT 50.486 69.756 67.408 69.845 ;
        RECT 50.44 69.802 67.362 69.891 ;
        RECT 50.394 69.848 67.316 69.937 ;
        RECT 50.348 69.894 67.27 69.983 ;
        RECT 50.302 69.94 67.224 70.029 ;
        RECT 50.256 69.986 67.178 70.075 ;
        RECT 50.21 70.032 67.132 70.121 ;
        RECT 50.164 70.078 67.086 70.167 ;
        RECT 50.118 70.124 67.04 70.213 ;
        RECT 50.072 70.17 66.994 70.259 ;
        RECT 50.026 70.216 66.948 70.305 ;
        RECT 49.98 70.262 66.902 70.351 ;
        RECT 49.934 70.308 66.856 70.397 ;
        RECT 49.888 70.354 66.81 70.443 ;
        RECT 49.842 70.4 66.764 70.489 ;
        RECT 49.796 70.446 66.718 70.535 ;
        RECT 49.75 70.492 66.672 70.581 ;
        RECT 49.704 70.538 66.626 70.627 ;
        RECT 49.658 70.584 66.58 70.673 ;
        RECT 49.612 70.63 66.534 70.719 ;
        RECT 49.566 70.676 66.488 70.765 ;
        RECT 49.52 70.722 66.442 70.811 ;
        RECT 49.474 70.768 66.396 70.857 ;
        RECT 49.428 70.814 66.35 70.903 ;
        RECT 49.382 70.86 66.304 70.949 ;
        RECT 49.336 70.906 66.258 70.995 ;
        RECT 49.29 70.952 66.212 71.041 ;
        RECT 49.244 70.998 66.166 71.087 ;
        RECT 49.198 71.044 66.12 71.133 ;
        RECT 49.152 71.09 66.074 71.179 ;
        RECT 49.106 71.136 66.028 71.225 ;
        RECT 49.06 71.182 65.982 71.271 ;
        RECT 49.014 71.228 65.936 71.317 ;
        RECT 48.968 71.274 65.89 71.363 ;
        RECT 48.922 71.32 65.844 71.409 ;
        RECT 48.876 71.366 65.798 71.455 ;
        RECT 48.83 71.412 65.752 71.501 ;
        RECT 48.784 71.458 65.706 71.547 ;
        RECT 48.738 71.504 65.66 71.593 ;
        RECT 48.692 71.55 65.614 71.639 ;
        RECT 48.646 71.596 65.568 71.685 ;
        RECT 48.6 71.642 65.522 71.731 ;
        RECT 48.554 71.688 65.476 71.777 ;
        RECT 48.508 71.734 65.43 71.823 ;
        RECT 48.462 71.78 65.384 71.869 ;
        RECT 48.416 71.826 65.338 71.915 ;
        RECT 48.37 71.872 65.292 71.961 ;
        RECT 48.324 71.918 65.246 72.007 ;
        RECT 48.278 71.964 65.2 72.053 ;
        RECT 48.232 72.01 65.154 72.099 ;
        RECT 48.186 72.056 65.108 72.145 ;
        RECT 48.14 72.102 65.062 72.191 ;
        RECT 48.094 72.148 65.016 72.237 ;
        RECT 48.048 72.194 64.97 72.283 ;
        RECT 48.002 72.24 64.924 72.329 ;
        RECT 47.956 72.286 64.878 72.375 ;
        RECT 47.91 72.332 64.832 72.421 ;
        RECT 47.864 72.378 64.786 72.467 ;
        RECT 47.818 72.424 64.74 72.513 ;
        RECT 47.772 72.47 64.694 72.559 ;
        RECT 47.726 72.516 64.648 72.605 ;
        RECT 47.68 72.562 64.602 72.651 ;
        RECT 47.634 72.608 64.556 72.697 ;
        RECT 47.588 72.654 64.51 72.743 ;
        RECT 47.542 72.7 64.464 72.789 ;
        RECT 47.496 72.746 64.418 72.835 ;
        RECT 47.45 72.792 64.372 72.881 ;
        RECT 47.404 72.838 64.326 72.927 ;
        RECT 47.358 72.884 64.28 72.973 ;
        RECT 47.312 72.93 64.234 73.019 ;
        RECT 47.266 72.976 64.188 73.065 ;
        RECT 47.22 73.022 64.142 73.111 ;
        RECT 47.174 73.068 64.096 73.157 ;
        RECT 47.128 73.114 64.05 73.203 ;
        RECT 47.082 73.16 64.004 73.249 ;
        RECT 47.036 73.206 63.958 73.295 ;
        RECT 46.99 73.252 63.912 73.341 ;
        RECT 46.944 73.298 63.866 73.387 ;
        RECT 46.898 73.344 63.82 73.433 ;
        RECT 46.852 73.39 63.774 73.479 ;
        RECT 46.806 73.436 63.728 73.525 ;
        RECT 46.76 73.482 63.682 73.571 ;
        RECT 46.714 73.528 63.636 73.617 ;
        RECT 46.668 73.574 63.59 73.663 ;
        RECT 46.622 73.62 63.544 73.709 ;
        RECT 46.576 73.666 63.498 73.755 ;
        RECT 46.53 73.712 63.452 73.801 ;
        RECT 46.484 73.758 63.406 73.847 ;
        RECT 46.438 73.804 63.36 73.893 ;
        RECT 46.392 73.85 63.314 73.939 ;
        RECT 46.346 73.896 63.268 73.985 ;
        RECT 46.3 73.942 63.222 74.031 ;
        RECT 46.254 73.988 63.176 74.077 ;
        RECT 46.208 74.034 63.13 74.123 ;
        RECT 46.162 74.08 63.084 74.169 ;
        RECT 46.116 74.126 63.038 74.215 ;
        RECT 46.07 74.172 62.992 74.261 ;
        RECT 46.024 74.218 62.946 74.307 ;
        RECT 45.978 74.264 62.9 74.353 ;
        RECT 45.932 74.31 62.854 74.399 ;
        RECT 45.886 74.356 62.808 74.445 ;
        RECT 45.84 74.402 62.762 74.491 ;
        RECT 45.794 74.448 62.716 74.537 ;
        RECT 45.748 74.494 62.67 74.583 ;
        RECT 45.702 74.54 62.624 74.629 ;
        RECT 45.656 74.586 62.578 74.675 ;
        RECT 45.61 74.632 62.532 74.721 ;
        RECT 45.564 74.678 62.486 74.767 ;
        RECT 45.518 74.724 62.44 74.813 ;
        RECT 45.472 74.77 62.394 74.859 ;
        RECT 45.426 74.816 62.348 74.905 ;
        RECT 45.38 74.862 62.302 74.951 ;
        RECT 45.334 74.908 62.256 74.997 ;
        RECT 45.288 74.954 62.21 75.043 ;
        RECT 45.242 75 62.164 75.089 ;
        RECT 45.196 75.046 62.118 75.135 ;
        RECT 45.15 75.092 62.072 75.181 ;
        RECT 45.104 75.138 62.026 75.227 ;
        RECT 45.058 75.184 61.98 75.273 ;
        RECT 45.012 75.23 61.934 75.319 ;
        RECT 44.966 75.276 61.888 75.365 ;
        RECT 44.92 75.322 61.842 75.411 ;
        RECT 44.874 75.368 61.796 75.457 ;
        RECT 44.828 75.414 61.75 75.503 ;
        RECT 44.782 75.46 61.704 75.549 ;
        RECT 44.736 75.506 61.658 75.595 ;
        RECT 44.69 75.552 61.612 75.641 ;
        RECT 44.644 75.598 61.566 75.687 ;
        RECT 44.598 75.644 61.52 75.733 ;
        RECT 44.552 75.69 61.474 75.779 ;
        RECT 44.506 75.736 61.428 75.825 ;
        RECT 44.46 75.782 61.382 75.871 ;
        RECT 44.414 75.828 61.336 75.917 ;
        RECT 44.368 75.874 61.29 75.963 ;
        RECT 44.322 75.92 61.244 76.009 ;
        RECT 44.276 75.966 61.198 76.055 ;
        RECT 44.23 76.012 61.152 76.101 ;
        RECT 44.184 76.058 61.106 76.147 ;
        RECT 44.138 76.104 61.06 76.193 ;
        RECT 44.092 76.15 61.014 76.239 ;
        RECT 44.046 76.196 60.968 76.285 ;
        RECT 44 76.242 60.922 76.331 ;
        RECT 44 76.242 60.876 76.377 ;
        RECT 44 76.242 60.83 76.423 ;
        RECT 44 76.242 60.784 76.469 ;
        RECT 44 76.242 60.738 76.515 ;
        RECT 44 76.242 60.692 76.561 ;
        RECT 44 76.242 60.646 76.607 ;
        RECT 44 76.242 60.6 76.653 ;
        RECT 44 76.242 60.554 76.699 ;
        RECT 44 76.242 60.508 76.745 ;
        RECT 44 76.242 60.462 76.791 ;
        RECT 44 76.242 60.416 76.837 ;
        RECT 44 76.242 60.37 76.883 ;
        RECT 44 76.242 60.324 76.929 ;
        RECT 44 76.242 60.278 76.975 ;
        RECT 44 76.242 60.232 77.021 ;
        RECT 44 76.242 60.186 77.067 ;
        RECT 44 76.242 60.14 77.113 ;
        RECT 44 76.242 60.094 77.159 ;
        RECT 44 76.242 60.048 77.205 ;
        RECT 44 76.242 60.002 77.251 ;
        RECT 44 76.242 59.956 77.297 ;
        RECT 44 76.242 59.91 77.343 ;
        RECT 44 76.242 59.864 77.389 ;
        RECT 44 76.242 59.818 77.435 ;
        RECT 44 76.242 59.772 77.481 ;
        RECT 44 76.242 59.726 77.527 ;
        RECT 44 76.242 59.68 77.573 ;
        RECT 44 76.242 59.634 77.619 ;
        RECT 44 76.242 59.588 77.665 ;
        RECT 44 76.242 59.542 77.711 ;
        RECT 44 76.242 59.496 77.757 ;
        RECT 44 76.242 59.45 77.803 ;
        RECT 44 76.242 59.404 77.849 ;
        RECT 44 76.242 59.358 77.895 ;
        RECT 44 76.242 59.312 77.941 ;
        RECT 44 76.242 59.266 77.987 ;
        RECT 44 76.242 59.22 78.033 ;
        RECT 44 76.242 59.174 78.079 ;
        RECT 44 76.242 59.128 78.125 ;
        RECT 44 76.242 59.082 78.171 ;
        RECT 44 76.242 59.036 78.217 ;
        RECT 44 76.242 58.99 78.263 ;
        RECT 44 76.242 58.944 78.309 ;
        RECT 44 76.242 58.898 78.355 ;
        RECT 44 76.242 58.852 78.401 ;
        RECT 44 76.242 58.806 78.447 ;
        RECT 44 76.242 58.76 78.493 ;
        RECT 44 76.242 58.714 78.539 ;
        RECT 44 76.242 58.668 78.585 ;
        RECT 44 76.242 58.622 78.631 ;
        RECT 44 76.242 58.576 78.677 ;
        RECT 44 76.242 58.53 78.723 ;
        RECT 44 76.242 58.484 78.769 ;
        RECT 44 76.242 58.438 78.815 ;
        RECT 44 76.242 58.392 78.861 ;
        RECT 44 76.242 58.346 78.907 ;
        RECT 44 76.242 58.3 78.953 ;
        RECT 44 76.242 58.254 78.999 ;
        RECT 44 76.242 58.208 79.045 ;
        RECT 44 76.242 58.162 79.091 ;
        RECT 44 76.242 58.116 79.137 ;
        RECT 44 76.242 58.07 79.183 ;
        RECT 44 76.242 58.024 79.229 ;
        RECT 44 76.242 57.978 79.275 ;
        RECT 44 76.242 57.932 79.321 ;
        RECT 44 76.242 57.886 79.367 ;
        RECT 44 76.242 57.84 79.413 ;
        RECT 44 76.242 57.794 79.459 ;
        RECT 44 76.242 57.748 79.505 ;
        RECT 44 76.242 57.702 79.551 ;
        RECT 44 76.242 57.656 79.597 ;
        RECT 44 76.242 57.61 79.643 ;
        RECT 44 76.242 57.564 79.689 ;
        RECT 44 76.242 57.518 79.735 ;
        RECT 44 76.242 57.472 79.781 ;
        RECT 44 76.242 57.426 79.827 ;
        RECT 44 76.242 57.38 79.873 ;
        RECT 44 76.242 57.334 79.919 ;
        RECT 44 76.242 57.288 79.965 ;
        RECT 44 76.242 57.242 80.011 ;
        RECT 44 76.242 57.196 80.057 ;
        RECT 44 76.242 57.15 80.103 ;
        RECT 44 76.242 57.104 80.149 ;
        RECT 44 76.242 57.058 80.195 ;
        RECT 44 76.242 57.012 80.241 ;
        RECT 44 76.242 56.966 80.287 ;
        RECT 44 76.242 56.92 80.333 ;
        RECT 44 76.242 56.874 80.379 ;
        RECT 44 76.242 56.828 80.425 ;
        RECT 44 76.242 56.782 80.471 ;
        RECT 44 76.242 56.736 80.517 ;
        RECT 44 76.242 56.69 80.563 ;
        RECT 44 76.242 56.644 80.609 ;
        RECT 44 76.242 56.598 80.655 ;
        RECT 44 76.242 56.552 80.701 ;
        RECT 44 76.242 56.506 80.747 ;
        RECT 44 76.242 56.46 80.793 ;
        RECT 44 76.242 56.414 80.839 ;
        RECT 44 76.242 56.368 80.885 ;
        RECT 44 76.242 56.322 80.931 ;
        RECT 44 76.242 56.276 80.977 ;
        RECT 44 76.242 56.23 81.023 ;
        RECT 44 76.242 56.184 81.069 ;
        RECT 44 76.242 56.138 81.115 ;
        RECT 44 76.242 56.092 81.161 ;
        RECT 44 76.242 56.046 81.207 ;
        RECT 44 76.242 56 110 ;
        RECT 82.76 57.5 110 63.5 ;
        RECT 76.748 63.489 85.24 63.521 ;
        RECT 74.31 65.927 82.76 65.996 ;
        RECT 74.356 65.881 82.806 65.957 ;
        RECT 82.728 57.516 82.76 65.996 ;
        RECT 74.264 65.973 82.728 66.035 ;
        RECT 74.402 65.835 82.852 65.911 ;
        RECT 82.682 57.555 82.728 66.035 ;
        RECT 74.218 66.019 82.682 66.081 ;
        RECT 74.448 65.789 82.898 65.865 ;
        RECT 82.636 57.601 82.682 66.081 ;
        RECT 74.172 66.065 82.636 66.127 ;
        RECT 74.494 65.743 82.944 65.819 ;
        RECT 82.59 57.647 82.636 66.127 ;
        RECT 74.126 66.111 82.59 66.173 ;
        RECT 74.54 65.697 82.99 65.773 ;
        RECT 82.544 57.693 82.59 66.173 ;
        RECT 74.08 66.157 82.544 66.219 ;
        RECT 74.586 65.651 83.036 65.727 ;
        RECT 82.498 57.739 82.544 66.219 ;
        RECT 74.034 66.203 82.498 66.265 ;
        RECT 74.632 65.605 83.082 65.681 ;
        RECT 82.452 57.785 82.498 66.265 ;
        RECT 73.988 66.249 82.452 66.311 ;
        RECT 74.678 65.559 83.128 65.635 ;
        RECT 82.406 57.831 82.452 66.311 ;
        RECT 73.942 66.295 82.406 66.357 ;
        RECT 74.724 65.513 83.174 65.589 ;
        RECT 82.36 57.877 82.406 66.357 ;
        RECT 73.896 66.341 82.36 66.403 ;
        RECT 74.77 65.467 83.22 65.543 ;
        RECT 82.314 57.923 82.36 66.403 ;
        RECT 73.85 66.387 82.314 66.449 ;
        RECT 74.816 65.421 83.266 65.497 ;
        RECT 82.268 57.969 82.314 66.449 ;
        RECT 73.804 66.433 82.268 66.495 ;
        RECT 74.862 65.375 83.312 65.451 ;
        RECT 82.222 58.015 82.268 66.495 ;
        RECT 73.758 66.479 82.222 66.541 ;
        RECT 74.908 65.329 83.358 65.405 ;
        RECT 82.176 58.061 82.222 66.541 ;
        RECT 73.712 66.525 82.176 66.587 ;
        RECT 74.954 65.283 83.404 65.359 ;
        RECT 82.13 58.107 82.176 66.587 ;
        RECT 73.666 66.571 82.13 66.633 ;
        RECT 75 65.237 83.45 65.313 ;
        RECT 82.084 58.153 82.13 66.633 ;
        RECT 73.62 66.617 82.084 66.679 ;
        RECT 75.046 65.191 83.496 65.267 ;
        RECT 82.038 58.199 82.084 66.679 ;
        RECT 73.574 66.663 82.038 66.725 ;
        RECT 75.092 65.145 83.542 65.221 ;
        RECT 81.992 58.245 82.038 66.725 ;
        RECT 73.528 66.709 81.992 66.771 ;
        RECT 75.138 65.099 83.588 65.175 ;
        RECT 81.946 58.291 81.992 66.771 ;
        RECT 73.482 66.755 81.946 66.817 ;
        RECT 75.184 65.053 83.634 65.129 ;
        RECT 81.9 58.337 81.946 66.817 ;
        RECT 73.436 66.801 81.9 66.863 ;
        RECT 75.23 65.007 83.68 65.083 ;
        RECT 81.854 58.383 81.9 66.863 ;
        RECT 73.39 66.847 81.854 66.909 ;
        RECT 75.276 64.961 83.726 65.037 ;
        RECT 81.808 58.429 81.854 66.909 ;
        RECT 73.344 66.893 81.808 66.955 ;
        RECT 75.322 64.915 83.772 64.991 ;
        RECT 81.762 58.475 81.808 66.955 ;
        RECT 73.298 66.939 81.762 67.001 ;
        RECT 75.368 64.869 83.818 64.945 ;
        RECT 81.716 58.521 81.762 67.001 ;
        RECT 73.252 66.985 81.716 67.047 ;
        RECT 75.414 64.823 83.864 64.899 ;
        RECT 81.67 58.567 81.716 67.047 ;
        RECT 73.206 67.031 81.67 67.093 ;
        RECT 75.46 64.777 83.91 64.853 ;
        RECT 81.624 58.613 81.67 67.093 ;
        RECT 73.16 67.077 81.624 67.139 ;
        RECT 75.506 64.731 83.956 64.807 ;
        RECT 81.578 58.659 81.624 67.139 ;
        RECT 73.114 67.123 81.578 67.185 ;
        RECT 75.552 64.685 84.002 64.761 ;
        RECT 81.532 58.705 81.578 67.185 ;
        RECT 73.068 67.169 81.532 67.231 ;
        RECT 75.598 64.639 84.048 64.715 ;
        RECT 81.486 58.751 81.532 67.231 ;
        RECT 73.022 67.215 81.486 67.277 ;
        RECT 75.644 64.593 84.094 64.669 ;
        RECT 81.44 58.797 81.486 67.277 ;
        RECT 72.976 67.261 81.44 67.323 ;
        RECT 75.69 64.547 84.14 64.623 ;
        RECT 81.394 58.843 81.44 67.323 ;
        RECT 72.93 67.307 81.394 67.369 ;
        RECT 75.736 64.501 84.186 64.577 ;
        RECT 81.348 58.889 81.394 67.369 ;
        RECT 72.884 67.353 81.348 67.415 ;
        RECT 75.782 64.455 84.232 64.531 ;
        RECT 81.302 58.935 81.348 67.415 ;
        RECT 72.838 67.399 81.302 67.461 ;
        RECT 75.828 64.409 84.278 64.485 ;
        RECT 81.256 58.981 81.302 67.461 ;
        RECT 72.792 67.445 81.256 67.507 ;
        RECT 75.874 64.363 84.324 64.439 ;
        RECT 81.21 59.027 81.256 67.507 ;
        RECT 72.746 67.491 81.21 67.553 ;
        RECT 75.92 64.317 84.37 64.393 ;
        RECT 81.164 59.073 81.21 67.553 ;
        RECT 72.7 67.537 81.164 67.599 ;
        RECT 75.966 64.271 84.416 64.347 ;
        RECT 81.118 59.119 81.164 67.599 ;
        RECT 72.654 67.583 81.118 67.645 ;
        RECT 76.012 64.225 84.462 64.301 ;
        RECT 81.072 59.165 81.118 67.645 ;
        RECT 72.608 67.629 81.072 67.691 ;
        RECT 76.058 64.179 84.508 64.255 ;
        RECT 81.026 59.211 81.072 67.691 ;
        RECT 72.562 67.675 81.026 67.737 ;
        RECT 76.104 64.133 84.554 64.209 ;
        RECT 80.98 59.257 81.026 67.737 ;
        RECT 72.516 67.721 80.98 67.783 ;
        RECT 76.15 64.087 84.6 64.163 ;
        RECT 80.934 59.303 80.98 67.783 ;
        RECT 72.47 67.767 80.934 67.829 ;
        RECT 76.196 64.041 84.646 64.117 ;
        RECT 80.888 59.349 80.934 67.829 ;
        RECT 72.424 67.813 80.888 67.875 ;
        RECT 76.242 63.995 84.692 64.071 ;
        RECT 80.842 59.395 80.888 67.875 ;
        RECT 72.378 67.859 80.842 67.921 ;
        RECT 76.288 63.949 84.738 64.025 ;
        RECT 80.796 59.441 80.842 67.921 ;
        RECT 72.332 67.905 80.796 67.967 ;
        RECT 76.334 63.903 84.784 63.979 ;
        RECT 80.75 59.487 80.796 67.967 ;
        RECT 72.286 67.951 80.75 68.013 ;
        RECT 76.38 63.857 84.83 63.933 ;
        RECT 80.704 59.533 80.75 68.013 ;
        RECT 72.24 67.997 80.704 68.059 ;
        RECT 76.426 63.811 84.876 63.887 ;
        RECT 80.658 59.579 80.704 68.059 ;
        RECT 72.194 68.043 80.658 68.105 ;
        RECT 76.472 63.765 84.922 63.841 ;
        RECT 80.612 59.625 80.658 68.105 ;
        RECT 72.148 68.089 80.612 68.151 ;
        RECT 76.518 63.719 84.968 63.795 ;
        RECT 80.566 59.671 80.612 68.151 ;
        RECT 72.102 68.135 80.566 68.197 ;
        RECT 76.564 63.673 85.014 63.749 ;
        RECT 80.52 59.717 80.566 68.197 ;
        RECT 72.056 68.181 80.52 68.243 ;
        RECT 76.61 63.627 85.06 63.703 ;
        RECT 80.474 59.763 80.52 68.243 ;
        RECT 72.01 68.227 80.474 68.289 ;
        RECT 76.656 63.581 85.106 63.657 ;
        RECT 80.428 59.809 80.474 68.289 ;
        RECT 71.964 68.273 80.428 68.335 ;
        RECT 76.702 63.535 85.152 63.611 ;
        RECT 80.382 59.855 80.428 68.335 ;
        RECT 71.918 68.319 80.382 68.381 ;
        RECT 76.748 63.489 85.198 63.565 ;
        RECT 80.336 59.901 80.382 68.381 ;
        RECT 71.872 68.365 80.336 68.427 ;
        RECT 76.794 63.443 110 63.5 ;
        RECT 80.29 59.947 80.336 68.427 ;
        RECT 71.826 68.411 80.29 68.473 ;
        RECT 76.84 63.397 110 63.5 ;
        RECT 80.244 59.993 80.29 68.473 ;
        RECT 71.78 68.457 80.244 68.519 ;
        RECT 76.886 63.351 110 63.5 ;
        RECT 80.198 60.039 80.244 68.519 ;
        RECT 71.734 68.503 80.198 68.565 ;
        RECT 76.932 63.305 110 63.5 ;
        RECT 80.152 60.085 80.198 68.565 ;
        RECT 71.688 68.549 80.152 68.611 ;
        RECT 76.978 63.259 110 63.5 ;
        RECT 80.106 60.131 80.152 68.611 ;
        RECT 71.642 68.595 80.106 68.657 ;
        RECT 77.024 63.213 110 63.5 ;
        RECT 80.06 60.177 80.106 68.657 ;
        RECT 71.596 68.641 80.06 68.703 ;
        RECT 77.07 63.167 110 63.5 ;
        RECT 80.014 60.223 80.06 68.703 ;
        RECT 71.55 68.687 80.014 68.749 ;
        RECT 77.116 63.121 110 63.5 ;
        RECT 79.968 60.269 80.014 68.749 ;
        RECT 71.504 68.733 79.968 68.795 ;
        RECT 77.162 63.075 110 63.5 ;
        RECT 79.922 60.315 79.968 68.795 ;
        RECT 71.458 68.779 79.922 68.841 ;
        RECT 77.208 63.029 110 63.5 ;
        RECT 79.876 60.361 79.922 68.841 ;
        RECT 71.412 68.825 79.876 68.887 ;
        RECT 77.254 62.983 110 63.5 ;
        RECT 79.83 60.407 79.876 68.887 ;
        RECT 71.366 68.871 79.83 68.933 ;
        RECT 77.3 62.937 110 63.5 ;
        RECT 79.784 60.453 79.83 68.933 ;
        RECT 71.32 68.917 79.784 68.979 ;
        RECT 77.346 62.891 110 63.5 ;
        RECT 79.738 60.499 79.784 68.979 ;
        RECT 71.274 68.963 79.738 69.025 ;
        RECT 77.392 62.845 110 63.5 ;
        RECT 79.692 60.545 79.738 69.025 ;
        RECT 71.228 69.009 79.692 69.071 ;
        RECT 77.438 62.799 110 63.5 ;
        RECT 79.646 60.591 79.692 69.071 ;
        RECT 71.182 69.055 79.646 69.117 ;
        RECT 77.484 62.753 110 63.5 ;
        RECT 79.6 60.637 79.646 69.117 ;
        RECT 71.136 69.101 79.6 69.163 ;
        RECT 77.53 62.707 110 63.5 ;
        RECT 79.554 60.683 79.6 69.163 ;
        RECT 71.09 69.147 79.554 69.209 ;
        RECT 77.576 62.661 110 63.5 ;
        RECT 79.508 60.729 79.554 69.209 ;
        RECT 71.044 69.193 79.508 69.255 ;
        RECT 77.622 62.615 110 63.5 ;
        RECT 79.462 60.775 79.508 69.255 ;
        RECT 70.998 69.239 79.462 69.301 ;
        RECT 77.668 62.569 110 63.5 ;
        RECT 79.416 60.821 79.462 69.301 ;
        RECT 70.952 69.285 79.416 69.347 ;
        RECT 77.714 62.523 110 63.5 ;
        RECT 79.37 60.867 79.416 69.347 ;
        RECT 70.906 69.331 79.37 69.393 ;
        RECT 77.76 62.477 110 63.5 ;
        RECT 79.324 60.913 79.37 69.393 ;
        RECT 70.86 69.377 79.324 69.439 ;
        RECT 77.806 62.431 110 63.5 ;
        RECT 79.278 60.959 79.324 69.439 ;
        RECT 70.814 69.423 79.278 69.485 ;
        RECT 77.852 62.385 110 63.5 ;
        RECT 69.515 30.5 110 42.5 ;
        RECT 57.496 42.496 74.48 42.522 ;
        RECT 52.574 47.418 69.515 47.472 ;
        RECT 52.62 47.372 69.561 47.442 ;
        RECT 69.502 30.506 69.515 47.472 ;
        RECT 52.666 47.326 69.607 47.396 ;
        RECT 69.456 30.536 69.502 47.501 ;
        RECT 52.528 47.464 69.456 47.547 ;
        RECT 52.712 47.28 69.653 47.35 ;
        RECT 69.41 30.582 69.456 47.547 ;
        RECT 52.482 47.51 69.41 47.593 ;
        RECT 52.758 47.234 69.699 47.304 ;
        RECT 69.364 30.628 69.41 47.593 ;
        RECT 52.436 47.556 69.364 47.639 ;
        RECT 52.804 47.188 69.745 47.258 ;
        RECT 69.318 30.674 69.364 47.639 ;
        RECT 52.39 47.602 69.318 47.685 ;
        RECT 52.85 47.142 69.791 47.212 ;
        RECT 69.272 30.72 69.318 47.685 ;
        RECT 52.344 47.648 69.272 47.731 ;
        RECT 52.896 47.096 69.837 47.166 ;
        RECT 69.226 30.766 69.272 47.731 ;
        RECT 52.298 47.694 69.226 47.777 ;
        RECT 52.942 47.05 69.883 47.12 ;
        RECT 69.18 30.812 69.226 47.777 ;
        RECT 52.252 47.74 69.18 47.823 ;
        RECT 52.988 47.004 69.929 47.074 ;
        RECT 69.134 30.858 69.18 47.823 ;
        RECT 52.206 47.786 69.134 47.869 ;
        RECT 53.034 46.958 69.975 47.028 ;
        RECT 69.088 30.904 69.134 47.869 ;
        RECT 52.16 47.832 69.088 47.915 ;
        RECT 53.08 46.912 70.021 46.982 ;
        RECT 69.042 30.95 69.088 47.915 ;
        RECT 52.114 47.878 69.042 47.961 ;
        RECT 53.126 46.866 70.067 46.936 ;
        RECT 68.996 30.996 69.042 47.961 ;
        RECT 52.068 47.924 68.996 48.007 ;
        RECT 53.172 46.82 70.113 46.89 ;
        RECT 68.95 31.042 68.996 48.007 ;
        RECT 52.022 47.97 68.95 48.053 ;
        RECT 53.218 46.774 70.159 46.844 ;
        RECT 68.904 31.088 68.95 48.053 ;
        RECT 51.976 48.016 68.904 48.099 ;
        RECT 53.264 46.728 70.205 46.798 ;
        RECT 68.858 31.134 68.904 48.099 ;
        RECT 51.93 48.062 68.858 48.145 ;
        RECT 53.31 46.682 70.251 46.752 ;
        RECT 68.812 31.18 68.858 48.145 ;
        RECT 51.884 48.108 68.812 48.191 ;
        RECT 53.356 46.636 70.297 46.706 ;
        RECT 68.766 31.226 68.812 48.191 ;
        RECT 51.838 48.154 68.766 48.237 ;
        RECT 53.402 46.59 70.343 46.66 ;
        RECT 68.72 31.272 68.766 48.237 ;
        RECT 51.792 48.2 68.72 48.283 ;
        RECT 53.448 46.544 70.389 46.614 ;
        RECT 68.674 31.318 68.72 48.283 ;
        RECT 51.746 48.246 68.674 48.329 ;
        RECT 53.494 46.498 70.435 46.568 ;
        RECT 68.628 31.364 68.674 48.329 ;
        RECT 51.7 48.292 68.628 48.375 ;
        RECT 53.54 46.452 70.481 46.522 ;
        RECT 68.582 31.41 68.628 48.375 ;
        RECT 51.654 48.338 68.582 48.421 ;
        RECT 53.586 46.406 70.527 46.476 ;
        RECT 68.536 31.456 68.582 48.421 ;
        RECT 51.608 48.384 68.536 48.467 ;
        RECT 53.632 46.36 70.573 46.43 ;
        RECT 68.49 31.502 68.536 48.467 ;
        RECT 51.562 48.43 68.49 48.513 ;
        RECT 53.678 46.314 70.619 46.384 ;
        RECT 68.444 31.548 68.49 48.513 ;
        RECT 51.516 48.476 68.444 48.559 ;
        RECT 53.724 46.268 70.665 46.338 ;
        RECT 68.398 31.594 68.444 48.559 ;
        RECT 51.47 48.522 68.398 48.605 ;
        RECT 53.77 46.222 70.711 46.292 ;
        RECT 68.352 31.64 68.398 48.605 ;
        RECT 51.424 48.568 68.352 48.651 ;
        RECT 53.816 46.176 70.757 46.246 ;
        RECT 68.306 31.686 68.352 48.651 ;
        RECT 51.378 48.614 68.306 48.697 ;
        RECT 53.862 46.13 70.803 46.2 ;
        RECT 68.26 31.732 68.306 48.697 ;
        RECT 51.332 48.66 68.26 48.743 ;
        RECT 53.908 46.084 70.849 46.154 ;
        RECT 68.214 31.778 68.26 48.743 ;
        RECT 51.286 48.706 68.214 48.789 ;
        RECT 53.954 46.038 70.895 46.108 ;
        RECT 68.168 31.824 68.214 48.789 ;
        RECT 51.24 48.752 68.168 48.835 ;
        RECT 54 45.992 70.941 46.062 ;
        RECT 68.122 31.87 68.168 48.835 ;
        RECT 51.194 48.798 68.122 48.881 ;
        RECT 54.046 45.946 70.987 46.016 ;
        RECT 68.076 31.916 68.122 48.881 ;
        RECT 51.148 48.844 68.076 48.927 ;
        RECT 54.092 45.9 71.033 45.97 ;
        RECT 68.03 31.962 68.076 48.927 ;
        RECT 51.102 48.89 68.03 48.973 ;
        RECT 54.138 45.854 71.079 45.924 ;
        RECT 67.984 32.008 68.03 48.973 ;
        RECT 51.056 48.936 67.984 49.019 ;
        RECT 54.184 45.808 71.125 45.878 ;
        RECT 67.938 32.054 67.984 49.019 ;
        RECT 51.01 48.982 67.938 49.065 ;
        RECT 54.23 45.762 71.171 45.832 ;
        RECT 67.892 32.1 67.938 49.065 ;
        RECT 50.964 49.028 67.892 49.111 ;
        RECT 54.276 45.716 71.217 45.786 ;
        RECT 67.846 32.146 67.892 49.111 ;
        RECT 50.918 49.074 67.846 49.157 ;
        RECT 54.322 45.67 71.263 45.74 ;
        RECT 67.8 32.192 67.846 49.157 ;
        RECT 50.872 49.12 67.8 49.203 ;
        RECT 54.368 45.624 71.309 45.694 ;
        RECT 67.754 32.238 67.8 49.203 ;
        RECT 50.826 49.166 67.754 49.249 ;
        RECT 54.414 45.578 71.355 45.648 ;
        RECT 67.708 32.284 67.754 49.249 ;
        RECT 50.78 49.212 67.708 49.295 ;
        RECT 54.46 45.532 71.401 45.602 ;
        RECT 67.662 32.33 67.708 49.295 ;
        RECT 50.734 49.258 67.662 49.341 ;
        RECT 54.506 45.486 71.447 45.556 ;
        RECT 67.616 32.376 67.662 49.341 ;
        RECT 50.688 49.304 67.616 49.387 ;
        RECT 54.552 45.44 71.493 45.51 ;
        RECT 67.57 32.422 67.616 49.387 ;
        RECT 50.642 49.35 67.57 49.433 ;
        RECT 54.598 45.394 71.539 45.464 ;
        RECT 67.524 32.468 67.57 49.433 ;
        RECT 50.596 49.396 67.524 49.479 ;
        RECT 54.644 45.348 71.585 45.418 ;
        RECT 67.478 32.514 67.524 49.479 ;
        RECT 50.55 49.442 67.478 49.525 ;
        RECT 54.69 45.302 71.631 45.372 ;
        RECT 67.432 32.56 67.478 49.525 ;
        RECT 50.504 49.488 67.432 49.571 ;
        RECT 54.736 45.256 71.677 45.326 ;
        RECT 67.386 32.606 67.432 49.571 ;
        RECT 50.458 49.534 67.386 49.617 ;
        RECT 54.782 45.21 71.723 45.28 ;
        RECT 67.34 32.652 67.386 49.617 ;
        RECT 50.412 49.58 67.34 49.663 ;
        RECT 54.828 45.164 71.769 45.234 ;
        RECT 67.294 32.698 67.34 49.663 ;
        RECT 50.366 49.626 67.294 49.709 ;
        RECT 54.874 45.118 71.815 45.188 ;
        RECT 67.248 32.744 67.294 49.709 ;
        RECT 50.32 49.672 67.248 49.755 ;
        RECT 54.92 45.072 71.861 45.142 ;
        RECT 67.202 32.79 67.248 49.755 ;
        RECT 50.274 49.718 67.202 49.801 ;
        RECT 54.966 45.026 71.907 45.096 ;
        RECT 67.156 32.836 67.202 49.801 ;
        RECT 50.228 49.764 67.156 49.847 ;
        RECT 55.012 44.98 71.953 45.05 ;
        RECT 67.11 32.882 67.156 49.847 ;
        RECT 50.182 49.81 67.11 49.893 ;
        RECT 55.058 44.934 71.999 45.004 ;
        RECT 67.064 32.928 67.11 49.893 ;
        RECT 50.136 49.856 67.064 49.939 ;
        RECT 55.104 44.888 72.045 44.958 ;
        RECT 67.018 32.974 67.064 49.939 ;
        RECT 50.09 49.902 67.018 49.985 ;
        RECT 55.15 44.842 72.091 44.912 ;
        RECT 66.972 33.02 67.018 49.985 ;
        RECT 50.044 49.948 66.972 50.031 ;
        RECT 55.196 44.796 72.137 44.866 ;
        RECT 66.926 33.066 66.972 50.031 ;
        RECT 49.998 49.994 66.926 50.077 ;
        RECT 55.242 44.75 72.183 44.82 ;
        RECT 66.88 33.112 66.926 50.077 ;
        RECT 49.952 50.04 66.88 50.123 ;
        RECT 55.288 44.704 72.229 44.774 ;
        RECT 66.834 33.158 66.88 50.123 ;
        RECT 49.906 50.086 66.834 50.169 ;
        RECT 55.334 44.658 72.275 44.728 ;
        RECT 66.788 33.204 66.834 50.169 ;
        RECT 49.86 50.132 66.788 50.215 ;
        RECT 55.38 44.612 72.321 44.682 ;
        RECT 66.742 33.25 66.788 50.215 ;
        RECT 49.814 50.178 66.742 50.261 ;
        RECT 55.426 44.566 72.367 44.636 ;
        RECT 66.696 33.296 66.742 50.261 ;
        RECT 49.768 50.224 66.696 50.307 ;
        RECT 55.472 44.52 72.413 44.59 ;
        RECT 66.65 33.342 66.696 50.307 ;
        RECT 49.722 50.27 66.65 50.353 ;
        RECT 55.518 44.474 72.459 44.544 ;
        RECT 66.604 33.388 66.65 50.353 ;
        RECT 49.676 50.316 66.604 50.399 ;
        RECT 55.564 44.428 72.505 44.498 ;
        RECT 66.558 33.434 66.604 50.399 ;
        RECT 49.63 50.362 66.558 50.445 ;
        RECT 55.61 44.382 72.551 44.452 ;
        RECT 66.512 33.48 66.558 50.445 ;
        RECT 49.584 50.408 66.512 50.491 ;
        RECT 55.656 44.336 72.597 44.406 ;
        RECT 66.466 33.526 66.512 50.491 ;
        RECT 49.538 50.454 66.466 50.537 ;
        RECT 55.702 44.29 72.643 44.36 ;
        RECT 66.42 33.572 66.466 50.537 ;
        RECT 49.492 50.5 66.42 50.583 ;
        RECT 55.748 44.244 72.689 44.314 ;
        RECT 66.374 33.618 66.42 50.583 ;
        RECT 49.446 50.546 66.374 50.629 ;
        RECT 55.794 44.198 72.735 44.268 ;
        RECT 66.328 33.664 66.374 50.629 ;
        RECT 49.4 50.592 66.328 50.675 ;
        RECT 55.84 44.152 72.781 44.222 ;
        RECT 66.282 33.71 66.328 50.675 ;
        RECT 49.354 50.638 66.282 50.721 ;
        RECT 55.886 44.106 72.827 44.176 ;
        RECT 66.236 33.756 66.282 50.721 ;
        RECT 49.308 50.684 66.236 50.767 ;
        RECT 55.932 44.06 72.873 44.13 ;
        RECT 66.19 33.802 66.236 50.767 ;
        RECT 49.262 50.73 66.19 50.813 ;
        RECT 55.978 44.014 72.919 44.084 ;
        RECT 66.144 33.848 66.19 50.813 ;
        RECT 49.216 50.776 66.144 50.859 ;
        RECT 56.024 43.968 72.965 44.038 ;
        RECT 66.098 33.894 66.144 50.859 ;
        RECT 49.17 50.822 66.098 50.905 ;
        RECT 56.07 43.922 73.011 43.992 ;
        RECT 66.052 33.94 66.098 50.905 ;
        RECT 49.124 50.868 66.052 50.951 ;
        RECT 56.116 43.876 73.057 43.946 ;
        RECT 66.006 33.986 66.052 50.951 ;
        RECT 49.078 50.914 66.006 50.997 ;
        RECT 56.162 43.83 73.103 43.9 ;
        RECT 65.96 34.032 66.006 50.997 ;
        RECT 49.032 50.96 65.96 51.043 ;
        RECT 56.208 43.784 73.149 43.854 ;
        RECT 65.914 34.078 65.96 51.043 ;
        RECT 48.986 51.006 65.914 51.089 ;
        RECT 56.254 43.738 73.195 43.808 ;
        RECT 65.868 34.124 65.914 51.089 ;
        RECT 48.94 51.052 65.868 51.135 ;
        RECT 56.3 43.692 73.241 43.762 ;
        RECT 65.822 34.17 65.868 51.135 ;
        RECT 48.894 51.098 65.822 51.181 ;
        RECT 56.346 43.646 73.287 43.716 ;
        RECT 65.776 34.216 65.822 51.181 ;
        RECT 48.848 51.144 65.776 51.227 ;
        RECT 56.392 43.6 73.333 43.67 ;
        RECT 65.73 34.262 65.776 51.227 ;
        RECT 48.802 51.19 65.73 51.273 ;
        RECT 56.438 43.554 73.379 43.624 ;
        RECT 65.684 34.308 65.73 51.273 ;
        RECT 48.756 51.236 65.684 51.319 ;
        RECT 56.484 43.508 73.425 43.578 ;
        RECT 65.638 34.354 65.684 51.319 ;
        RECT 48.71 51.282 65.638 51.365 ;
        RECT 56.53 43.462 73.471 43.532 ;
        RECT 65.592 34.4 65.638 51.365 ;
        RECT 48.664 51.328 65.592 51.411 ;
        RECT 56.576 43.416 73.517 43.486 ;
        RECT 65.546 34.446 65.592 51.411 ;
        RECT 48.618 51.374 65.546 51.457 ;
        RECT 56.622 43.37 73.563 43.44 ;
        RECT 65.5 34.492 65.546 51.457 ;
        RECT 48.572 51.42 65.5 51.503 ;
        RECT 56.668 43.324 73.609 43.394 ;
        RECT 65.454 34.538 65.5 51.503 ;
        RECT 48.526 51.466 65.454 51.549 ;
        RECT 56.714 43.278 73.655 43.348 ;
        RECT 65.408 34.584 65.454 51.549 ;
        RECT 48.48 51.512 65.408 51.595 ;
        RECT 56.76 43.232 73.701 43.302 ;
        RECT 65.362 34.63 65.408 51.595 ;
        RECT 48.434 51.558 65.362 51.641 ;
        RECT 56.806 43.186 73.747 43.256 ;
        RECT 65.316 34.676 65.362 51.641 ;
        RECT 48.388 51.604 65.316 51.687 ;
        RECT 56.852 43.14 73.793 43.21 ;
        RECT 65.27 34.722 65.316 51.687 ;
        RECT 48.342 51.65 65.27 51.733 ;
        RECT 56.898 43.094 73.839 43.164 ;
        RECT 65.224 34.768 65.27 51.733 ;
        RECT 48.296 51.696 65.224 51.779 ;
        RECT 56.944 43.048 73.885 43.118 ;
        RECT 65.178 34.814 65.224 51.779 ;
        RECT 48.25 51.742 65.178 51.825 ;
        RECT 56.99 43.002 73.931 43.072 ;
        RECT 65.132 34.86 65.178 51.825 ;
        RECT 48.204 51.788 65.132 51.871 ;
        RECT 57.036 42.956 73.977 43.026 ;
        RECT 65.086 34.906 65.132 51.871 ;
        RECT 48.158 51.834 65.086 51.917 ;
        RECT 57.082 42.91 74.023 42.98 ;
        RECT 65.04 34.952 65.086 51.917 ;
        RECT 48.112 51.88 65.04 51.963 ;
        RECT 57.128 42.864 74.069 42.934 ;
        RECT 64.994 34.998 65.04 51.963 ;
        RECT 48.066 51.926 64.994 52.009 ;
        RECT 57.174 42.818 74.115 42.888 ;
        RECT 64.948 35.044 64.994 52.009 ;
        RECT 48.02 51.972 64.948 52.055 ;
        RECT 57.22 42.772 74.161 42.842 ;
        RECT 64.902 35.09 64.948 52.055 ;
        RECT 47.974 52.018 64.902 52.101 ;
        RECT 57.266 42.726 74.207 42.796 ;
        RECT 64.856 35.136 64.902 52.101 ;
        RECT 47.928 52.064 64.856 52.147 ;
        RECT 57.312 42.68 74.253 42.75 ;
        RECT 64.81 35.182 64.856 52.147 ;
        RECT 47.882 52.11 64.81 52.193 ;
        RECT 57.358 42.634 74.299 42.704 ;
        RECT 64.764 35.228 64.81 52.193 ;
        RECT 47.836 52.156 64.764 52.239 ;
        RECT 57.404 42.588 74.345 42.658 ;
        RECT 64.718 35.274 64.764 52.239 ;
        RECT 47.79 52.202 64.718 52.285 ;
        RECT 57.45 42.542 74.391 42.612 ;
        RECT 64.672 35.32 64.718 52.285 ;
        RECT 47.744 52.248 64.672 52.331 ;
        RECT 57.496 42.496 74.437 42.566 ;
        RECT 64.626 35.366 64.672 52.331 ;
        RECT 47.698 52.294 64.626 52.377 ;
        RECT 57.542 42.45 110 42.5 ;
        RECT 64.58 35.412 64.626 52.377 ;
        RECT 47.652 52.34 64.58 52.423 ;
        RECT 57.588 42.404 110 42.5 ;
        RECT 64.534 35.458 64.58 52.423 ;
        RECT 47.606 52.386 64.534 52.469 ;
        RECT 57.634 42.358 110 42.5 ;
        RECT 64.488 35.504 64.534 52.469 ;
        RECT 47.56 52.432 64.488 52.515 ;
        RECT 57.68 42.312 110 42.5 ;
        RECT 64.442 35.55 64.488 52.515 ;
        RECT 47.514 52.478 64.442 52.561 ;
        RECT 57.726 42.266 110 42.5 ;
        RECT 64.396 35.596 64.442 52.561 ;
        RECT 47.468 52.524 64.396 52.607 ;
        RECT 57.772 42.22 110 42.5 ;
        RECT 64.35 35.642 64.396 52.607 ;
        RECT 47.422 52.57 64.35 52.653 ;
        RECT 57.818 42.174 110 42.5 ;
        RECT 64.304 35.688 64.35 52.653 ;
        RECT 47.376 52.616 64.304 52.699 ;
        RECT 57.864 42.128 110 42.5 ;
        RECT 64.258 35.734 64.304 52.699 ;
        RECT 47.33 52.662 64.258 52.745 ;
        RECT 57.91 42.082 110 42.5 ;
        RECT 64.212 35.78 64.258 52.745 ;
        RECT 47.284 52.708 64.212 52.791 ;
        RECT 57.956 42.036 110 42.5 ;
        RECT 64.166 35.826 64.212 52.791 ;
        RECT 47.238 52.754 64.166 52.837 ;
        RECT 58.002 41.99 110 42.5 ;
        RECT 64.12 35.872 64.166 52.837 ;
        RECT 47.192 52.8 64.12 52.883 ;
        RECT 58.048 41.944 110 42.5 ;
        RECT 64.074 35.918 64.12 52.883 ;
        RECT 47.146 52.846 64.074 52.929 ;
        RECT 58.094 41.898 110 42.5 ;
        RECT 64.028 35.964 64.074 52.929 ;
        RECT 47.1 52.892 64.028 52.975 ;
        RECT 58.14 41.852 110 42.5 ;
        RECT 63.982 36.01 64.028 52.975 ;
        RECT 47.054 52.938 63.982 53.021 ;
        RECT 58.186 41.806 110 42.5 ;
        RECT 63.936 36.056 63.982 53.021 ;
        RECT 47.008 52.984 63.936 53.067 ;
        RECT 58.232 41.76 110 42.5 ;
        RECT 63.89 36.102 63.936 53.067 ;
        RECT 46.962 53.03 63.89 53.113 ;
        RECT 58.278 41.714 110 42.5 ;
        RECT 63.844 36.148 63.89 53.113 ;
        RECT 46.916 53.076 63.844 53.159 ;
        RECT 58.324 41.668 110 42.5 ;
        RECT 63.798 36.194 63.844 53.159 ;
        RECT 46.87 53.122 63.798 53.205 ;
        RECT 58.37 41.622 110 42.5 ;
        RECT 63.752 36.24 63.798 53.205 ;
        RECT 46.824 53.168 63.752 53.251 ;
        RECT 58.416 41.576 110 42.5 ;
        RECT 63.706 36.286 63.752 53.251 ;
        RECT 46.778 53.214 63.706 53.297 ;
        RECT 58.462 41.53 110 42.5 ;
        RECT 63.66 36.332 63.706 53.297 ;
        RECT 46.732 53.26 63.66 53.343 ;
        RECT 58.508 41.484 110 42.5 ;
        RECT 63.614 36.378 63.66 53.343 ;
        RECT 46.686 53.306 63.614 53.389 ;
        RECT 58.554 41.438 110 42.5 ;
        RECT 63.568 36.424 63.614 53.389 ;
        RECT 46.64 53.352 63.568 53.435 ;
        RECT 58.6 41.392 110 42.5 ;
        RECT 63.522 36.47 63.568 53.435 ;
        RECT 46.594 53.398 63.522 53.481 ;
        RECT 58.646 41.346 110 42.5 ;
        RECT 63.476 36.516 63.522 53.481 ;
        RECT 46.548 53.444 63.476 53.527 ;
        RECT 58.692 41.3 110 42.5 ;
        RECT 63.43 36.562 63.476 53.527 ;
        RECT 46.502 53.49 63.43 53.573 ;
        RECT 58.738 41.254 110 42.5 ;
        RECT 63.384 36.608 63.43 53.573 ;
        RECT 46.456 53.536 63.384 53.619 ;
        RECT 58.784 41.208 110 42.5 ;
        RECT 63.338 36.654 63.384 53.619 ;
        RECT 46.41 53.582 63.338 53.665 ;
        RECT 58.83 41.162 110 42.5 ;
        RECT 63.292 36.7 63.338 53.665 ;
        RECT 46.364 53.628 63.292 53.711 ;
        RECT 58.876 41.116 110 42.5 ;
        RECT 63.246 36.746 63.292 53.711 ;
        RECT 46.318 53.674 63.246 53.757 ;
        RECT 58.922 41.07 110 42.5 ;
        RECT 63.2 36.792 63.246 53.757 ;
        RECT 46.272 53.72 63.2 53.803 ;
        RECT 58.968 41.024 110 42.5 ;
        RECT 63.154 36.838 63.2 53.803 ;
        RECT 46.226 53.766 63.154 53.849 ;
        RECT 59.014 40.978 110 42.5 ;
        RECT 63.108 36.884 63.154 53.849 ;
        RECT 46.18 53.812 63.108 53.895 ;
        RECT 59.06 40.932 110 42.5 ;
        RECT 63.062 36.93 63.108 53.895 ;
        RECT 46.134 53.858 63.062 53.941 ;
        RECT 59.106 40.886 110 42.5 ;
        RECT 63.016 36.976 63.062 53.941 ;
        RECT 46.088 53.904 63.016 53.987 ;
        RECT 59.152 40.84 110 42.5 ;
        RECT 62.97 37.022 63.016 53.987 ;
        RECT 46.042 53.95 62.97 54.033 ;
        RECT 59.198 40.794 110 42.5 ;
        RECT 62.924 37.068 62.97 54.033 ;
        RECT 45.996 53.996 62.924 54.079 ;
        RECT 59.244 40.748 110 42.5 ;
        RECT 62.878 37.114 62.924 54.079 ;
        RECT 45.95 54.042 62.878 54.125 ;
        RECT 59.29 40.702 110 42.5 ;
        RECT 62.832 37.16 62.878 54.125 ;
        RECT 45.904 54.088 62.832 54.171 ;
        RECT 59.336 40.656 110 42.5 ;
        RECT 62.786 37.206 62.832 54.171 ;
        RECT 45.858 54.134 62.786 54.217 ;
        RECT 59.382 40.61 110 42.5 ;
        RECT 62.74 37.252 62.786 54.217 ;
        RECT 45.812 54.18 62.74 54.263 ;
        RECT 59.428 40.564 110 42.5 ;
        RECT 62.694 37.298 62.74 54.263 ;
        RECT 45.766 54.226 62.694 54.309 ;
        RECT 59.474 40.518 110 42.5 ;
        RECT 62.648 37.344 62.694 54.309 ;
        RECT 45.72 54.272 62.648 54.355 ;
        RECT 59.52 40.472 110 42.5 ;
        RECT 62.602 37.39 62.648 54.355 ;
        RECT 45.674 54.318 62.602 54.401 ;
        RECT 59.566 40.426 110 42.5 ;
        RECT 62.556 37.436 62.602 54.401 ;
        RECT 45.628 54.364 62.556 54.447 ;
        RECT 59.612 40.38 110 42.5 ;
        RECT 62.51 37.482 62.556 54.447 ;
        RECT 45.582 54.41 62.51 54.493 ;
        RECT 59.658 40.334 110 42.5 ;
        RECT 62.464 37.528 62.51 54.493 ;
        RECT 45.536 54.456 62.464 54.539 ;
        RECT 59.704 40.288 110 42.5 ;
        RECT 62.418 37.574 62.464 54.539 ;
        RECT 45.49 54.502 62.418 54.585 ;
        RECT 59.75 40.242 110 42.5 ;
        RECT 62.372 37.62 62.418 54.585 ;
        RECT 45.444 54.548 62.372 54.631 ;
        RECT 59.796 40.196 110 42.5 ;
        RECT 62.326 37.666 62.372 54.631 ;
        RECT 45.398 54.594 62.326 54.677 ;
        RECT 59.842 40.15 110 42.5 ;
        RECT 62.28 37.712 62.326 54.677 ;
        RECT 45.352 54.64 62.28 54.723 ;
        RECT 59.888 40.104 110 42.5 ;
        RECT 62.234 37.758 62.28 54.723 ;
        RECT 45.306 54.686 62.234 54.769 ;
        RECT 59.934 40.058 110 42.5 ;
        RECT 62.188 37.804 62.234 54.769 ;
        RECT 45.26 54.732 62.188 54.815 ;
        RECT 59.98 40.012 110 42.5 ;
        RECT 62.142 37.85 62.188 54.815 ;
        RECT 45.214 54.778 62.142 54.861 ;
        RECT 60.026 39.966 110 42.5 ;
        RECT 62.096 37.896 62.142 54.861 ;
        RECT 45.168 54.824 62.096 54.907 ;
        RECT 60.072 39.92 110 42.5 ;
        RECT 62.05 37.942 62.096 54.907 ;
        RECT 45.122 54.87 62.05 54.953 ;
        RECT 60.118 39.874 110 42.5 ;
        RECT 62.004 37.988 62.05 54.953 ;
        RECT 45.076 54.916 62.004 54.999 ;
        RECT 60.164 39.828 110 42.5 ;
        RECT 61.958 38.034 62.004 54.999 ;
        RECT 45.03 54.962 61.958 55.045 ;
        RECT 60.21 39.782 110 42.5 ;
        RECT 61.912 38.08 61.958 55.045 ;
        RECT 44.984 55.008 61.912 55.091 ;
        RECT 60.256 39.736 110 42.5 ;
        RECT 61.866 38.126 61.912 55.091 ;
        RECT 44.938 55.054 61.866 55.137 ;
        RECT 60.302 39.69 110 42.5 ;
        RECT 61.82 38.172 61.866 55.137 ;
        RECT 44.892 55.1 61.82 55.183 ;
        RECT 60.348 39.644 110 42.5 ;
        RECT 61.774 38.218 61.82 55.183 ;
        RECT 44.846 55.146 61.774 55.229 ;
        RECT 60.394 39.598 110 42.5 ;
        RECT 61.728 38.264 61.774 55.229 ;
        RECT 44.8 55.192 61.728 55.275 ;
        RECT 60.44 39.552 110 42.5 ;
        RECT 61.682 38.31 61.728 55.275 ;
        RECT 44.754 55.238 61.682 55.321 ;
        RECT 60.486 39.506 110 42.5 ;
        RECT 61.636 38.356 61.682 55.321 ;
        RECT 44.708 55.284 61.636 55.367 ;
        RECT 60.532 39.46 110 42.5 ;
        RECT 61.59 38.402 61.636 55.367 ;
        RECT 44.662 55.33 61.59 55.413 ;
        RECT 60.578 39.414 110 42.5 ;
        RECT 61.544 38.448 61.59 55.413 ;
        RECT 44.616 55.376 61.544 55.459 ;
        RECT 60.624 39.368 110 42.5 ;
        RECT 61.498 38.494 61.544 55.459 ;
        RECT 44.57 55.422 61.498 55.505 ;
        RECT 60.67 39.322 110 42.5 ;
        RECT 61.452 38.54 61.498 55.505 ;
        RECT 44.524 55.468 61.452 55.551 ;
        RECT 60.716 39.276 110 42.5 ;
        RECT 61.406 38.586 61.452 55.551 ;
        RECT 44.478 55.514 61.406 55.597 ;
        RECT 60.762 39.23 110 42.5 ;
        RECT 61.36 38.632 61.406 55.597 ;
        RECT 44.432 55.56 61.36 55.643 ;
        RECT 60.808 39.184 110 42.5 ;
        RECT 61.314 38.678 61.36 55.643 ;
        RECT 44.386 55.606 61.314 55.689 ;
        RECT 60.854 39.138 110 42.5 ;
        RECT 61.268 38.724 61.314 55.689 ;
        RECT 44.34 55.652 61.268 55.735 ;
        RECT 60.9 39.092 110 42.5 ;
        RECT 61.222 38.77 61.268 55.735 ;
        RECT 44.294 55.698 61.222 55.781 ;
        RECT 60.946 39.046 110 42.5 ;
        RECT 61.176 38.816 61.222 55.781 ;
        RECT 44.248 55.744 61.176 55.827 ;
        RECT 60.992 39 110 42.5 ;
        RECT 61.13 38.862 61.176 55.827 ;
        RECT 44.202 55.79 61.13 55.873 ;
        RECT 61.038 38.954 110 42.5 ;
        RECT 61.084 38.908 61.13 55.873 ;
        RECT 44.156 55.836 61.084 55.919 ;
        RECT 44.11 55.882 61.038 55.965 ;
        RECT 44.064 55.928 60.992 56.011 ;
        RECT 44.018 55.974 60.946 56.057 ;
        RECT 43.972 56.02 60.9 56.103 ;
        RECT 43.926 56.066 60.854 56.149 ;
        RECT 43.88 56.112 60.808 56.195 ;
        RECT 43.834 56.158 60.762 56.241 ;
        RECT 43.788 56.204 60.716 56.287 ;
        RECT 43.742 56.25 60.67 56.333 ;
        RECT 43.696 56.296 60.624 56.379 ;
        RECT 43.65 56.342 60.578 56.425 ;
        RECT 43.604 56.388 60.532 56.471 ;
        RECT 43.558 56.434 60.486 56.517 ;
        RECT 43.512 56.48 60.44 56.563 ;
        RECT 43.466 56.526 60.394 56.609 ;
        RECT 43.42 56.572 60.348 56.655 ;
        RECT 43.374 56.618 60.302 56.701 ;
        RECT 43.328 56.664 60.256 56.747 ;
        RECT 43.282 56.71 60.21 56.793 ;
        RECT 43.236 56.756 60.164 56.839 ;
        RECT 43.19 56.802 60.118 56.885 ;
        RECT 43.144 56.848 60.072 56.931 ;
        RECT 43.098 56.894 60.026 56.977 ;
        RECT 43.052 56.94 59.98 57.023 ;
        RECT 43.006 56.986 59.934 57.069 ;
        RECT 42.96 57.032 59.888 57.115 ;
        RECT 42.914 57.078 59.842 57.161 ;
        RECT 42.868 57.124 59.796 57.207 ;
        RECT 42.822 57.17 59.75 57.253 ;
        RECT 42.776 57.216 59.704 57.299 ;
        RECT 42.73 57.262 59.658 57.345 ;
        RECT 42.684 57.308 59.612 57.391 ;
        RECT 42.638 57.354 59.566 57.437 ;
        RECT 42.592 57.4 59.52 57.483 ;
        RECT 42.546 57.446 59.474 57.529 ;
        RECT 42.5 57.492 59.428 57.575 ;
        RECT 42.46 57.535 59.382 57.621 ;
        RECT 42.414 57.578 59.336 57.667 ;
        RECT 42.368 57.624 59.29 57.713 ;
        RECT 42.322 57.67 59.244 57.759 ;
        RECT 42.276 57.716 59.198 57.805 ;
        RECT 42.23 57.762 59.152 57.851 ;
        RECT 42.184 57.808 59.106 57.897 ;
        RECT 42.138 57.854 59.06 57.943 ;
        RECT 42.092 57.9 59.014 57.989 ;
        RECT 42.046 57.946 58.968 58.035 ;
        RECT 42 57.992 58.922 58.081 ;
        RECT 41.954 58.038 58.876 58.127 ;
        RECT 41.908 58.084 58.83 58.173 ;
        RECT 41.862 58.13 58.784 58.219 ;
        RECT 41.816 58.176 58.738 58.265 ;
        RECT 41.77 58.222 58.692 58.311 ;
        RECT 41.724 58.268 58.646 58.357 ;
        RECT 41.678 58.314 58.6 58.403 ;
        RECT 41.632 58.36 58.554 58.449 ;
        RECT 41.586 58.406 58.508 58.495 ;
        RECT 41.54 58.452 58.462 58.541 ;
        RECT 41.494 58.498 58.416 58.587 ;
        RECT 41.448 58.544 58.37 58.633 ;
        RECT 41.402 58.59 58.324 58.679 ;
        RECT 41.356 58.636 58.278 58.725 ;
        RECT 41.31 58.682 58.232 58.771 ;
        RECT 41.264 58.728 58.186 58.817 ;
        RECT 41.218 58.774 58.14 58.863 ;
        RECT 41.172 58.82 58.094 58.909 ;
        RECT 41.126 58.866 58.048 58.955 ;
        RECT 41.08 58.912 58.002 59.001 ;
        RECT 41.034 58.958 57.956 59.047 ;
        RECT 40.988 59.004 57.91 59.093 ;
        RECT 40.942 59.05 57.864 59.139 ;
        RECT 40.896 59.096 57.818 59.185 ;
        RECT 40.85 59.142 57.772 59.231 ;
        RECT 40.804 59.188 57.726 59.277 ;
        RECT 40.758 59.234 57.68 59.323 ;
        RECT 40.712 59.28 57.634 59.369 ;
        RECT 40.666 59.326 57.588 59.415 ;
        RECT 40.62 59.372 57.542 59.461 ;
        RECT 40.574 59.418 57.496 59.507 ;
        RECT 40.528 59.464 57.45 59.553 ;
        RECT 40.482 59.51 57.404 59.599 ;
        RECT 40.436 59.556 57.358 59.645 ;
        RECT 40.39 59.602 57.312 59.691 ;
        RECT 40.344 59.648 57.266 59.737 ;
        RECT 40.298 59.694 57.22 59.783 ;
        RECT 40.252 59.74 57.174 59.829 ;
        RECT 40.206 59.786 57.128 59.875 ;
        RECT 40.16 59.832 57.082 59.921 ;
        RECT 40.114 59.878 57.036 59.967 ;
        RECT 40.068 59.924 56.99 60.013 ;
        RECT 40.022 59.97 56.944 60.059 ;
        RECT 39.976 60.016 56.898 60.105 ;
        RECT 39.93 60.062 56.852 60.151 ;
        RECT 39.884 60.108 56.806 60.197 ;
        RECT 39.838 60.154 56.76 60.243 ;
        RECT 39.792 60.2 56.714 60.289 ;
        RECT 39.746 60.246 56.668 60.335 ;
        RECT 39.7 60.292 56.622 60.381 ;
        RECT 39.654 60.338 56.576 60.427 ;
        RECT 39.608 60.384 56.53 60.473 ;
        RECT 39.562 60.43 56.484 60.519 ;
        RECT 39.516 60.476 56.438 60.565 ;
        RECT 39.47 60.522 56.392 60.611 ;
        RECT 39.424 60.568 56.346 60.657 ;
        RECT 39.378 60.614 56.3 60.703 ;
        RECT 39.332 60.66 56.254 60.749 ;
        RECT 39.286 60.706 56.208 60.795 ;
        RECT 39.24 60.752 56.162 60.841 ;
        RECT 39.194 60.798 56.116 60.887 ;
        RECT 39.148 60.844 56.07 60.933 ;
        RECT 39.102 60.89 56.024 60.979 ;
        RECT 39.056 60.936 55.978 61.025 ;
        RECT 39.01 60.982 55.932 61.071 ;
        RECT 38.964 61.028 55.886 61.117 ;
        RECT 38.918 61.074 55.84 61.163 ;
        RECT 38.872 61.12 55.794 61.209 ;
        RECT 38.826 61.166 55.748 61.255 ;
        RECT 38.78 61.212 55.702 61.301 ;
        RECT 38.734 61.258 55.656 61.347 ;
        RECT 38.688 61.304 55.61 61.393 ;
        RECT 38.642 61.35 55.564 61.439 ;
        RECT 38.596 61.396 55.518 61.485 ;
        RECT 38.55 61.442 55.472 61.531 ;
        RECT 38.504 61.488 55.426 61.577 ;
        RECT 38.458 61.534 55.38 61.623 ;
        RECT 38.412 61.58 55.334 61.669 ;
        RECT 38.366 61.626 55.288 61.715 ;
        RECT 38.32 61.672 55.242 61.761 ;
        RECT 38.274 61.718 55.196 61.807 ;
        RECT 38.228 61.764 55.15 61.853 ;
        RECT 38.182 61.81 55.104 61.899 ;
        RECT 38.136 61.856 55.058 61.945 ;
        RECT 38.09 61.902 55.012 61.991 ;
        RECT 38.044 61.948 54.966 62.037 ;
        RECT 37.998 61.994 54.92 62.083 ;
        RECT 37.952 62.04 54.874 62.129 ;
        RECT 37.906 62.086 54.828 62.175 ;
        RECT 37.86 62.132 54.782 62.221 ;
        RECT 37.814 62.178 54.736 62.267 ;
        RECT 37.768 62.224 54.69 62.313 ;
        RECT 37.722 62.27 54.644 62.359 ;
        RECT 37.676 62.316 54.598 62.405 ;
        RECT 37.63 62.362 54.552 62.451 ;
        RECT 37.584 62.408 54.506 62.497 ;
        RECT 37.538 62.454 54.46 62.543 ;
        RECT 37.492 62.5 54.414 62.589 ;
        RECT 37.446 62.546 54.368 62.635 ;
        RECT 37.4 62.592 54.322 62.681 ;
        RECT 37.354 62.638 54.276 62.727 ;
        RECT 37.308 62.684 54.23 62.773 ;
        RECT 37.262 62.73 54.184 62.819 ;
        RECT 37.216 62.776 54.138 62.865 ;
        RECT 37.17 62.822 54.092 62.911 ;
        RECT 37.124 62.868 54.046 62.957 ;
        RECT 37.078 62.914 54 63.003 ;
        RECT 37.032 62.96 53.954 63.049 ;
        RECT 36.986 63.006 53.908 63.095 ;
        RECT 36.94 63.052 53.862 63.141 ;
        RECT 36.894 63.098 53.816 63.187 ;
        RECT 36.848 63.144 53.77 63.233 ;
        RECT 36.802 63.19 53.724 63.279 ;
        RECT 36.756 63.236 53.678 63.325 ;
        RECT 36.71 63.282 53.632 63.371 ;
        RECT 36.664 63.328 53.586 63.417 ;
        RECT 36.618 63.374 53.54 63.463 ;
        RECT 36.572 63.42 53.494 63.509 ;
        RECT 36.526 63.466 53.448 63.555 ;
        RECT 36.48 63.512 53.402 63.601 ;
        RECT 36.434 63.558 53.356 63.647 ;
        RECT 36.388 63.604 53.31 63.693 ;
        RECT 36.342 63.65 53.264 63.739 ;
        RECT 36.296 63.696 53.218 63.785 ;
        RECT 36.25 63.742 53.172 63.831 ;
        RECT 36.204 63.788 53.126 63.877 ;
        RECT 36.158 63.834 53.08 63.923 ;
        RECT 36.112 63.88 53.034 63.969 ;
        RECT 36.066 63.926 52.988 64.015 ;
        RECT 36.02 63.972 52.942 64.061 ;
        RECT 35.974 64.018 52.896 64.107 ;
        RECT 35.928 64.064 52.85 64.153 ;
        RECT 35.882 64.11 52.804 64.199 ;
        RECT 35.836 64.156 52.758 64.245 ;
        RECT 35.79 64.202 52.712 64.291 ;
        RECT 35.744 64.248 52.666 64.337 ;
        RECT 35.698 64.294 52.62 64.383 ;
        RECT 35.652 64.34 52.574 64.429 ;
        RECT 35.606 64.386 52.528 64.475 ;
        RECT 35.56 64.432 52.482 64.521 ;
        RECT 35.514 64.478 52.436 64.567 ;
        RECT 35.468 64.524 52.39 64.613 ;
        RECT 35.422 64.57 52.344 64.659 ;
        RECT 35.376 64.616 52.298 64.705 ;
        RECT 35.33 64.662 52.252 64.751 ;
        RECT 35.284 64.708 52.206 64.797 ;
        RECT 35.238 64.754 52.16 64.843 ;
        RECT 35.192 64.8 52.114 64.889 ;
        RECT 35.146 64.846 52.068 64.935 ;
        RECT 35.1 64.892 52.022 64.981 ;
        RECT 35.054 64.938 51.976 65.027 ;
        RECT 35.008 64.984 51.93 65.073 ;
        RECT 34.962 65.03 51.884 65.119 ;
        RECT 34.916 65.076 51.838 65.165 ;
        RECT 34.87 65.122 51.792 65.211 ;
        RECT 34.824 65.168 51.746 65.257 ;
        RECT 34.778 65.214 51.7 65.303 ;
        RECT 34.732 65.26 51.654 65.349 ;
        RECT 34.686 65.306 51.608 65.395 ;
        RECT 34.64 65.352 51.562 65.441 ;
        RECT 34.594 65.398 51.516 65.487 ;
        RECT 34.548 65.444 51.47 65.533 ;
        RECT 34.502 65.49 51.424 65.579 ;
        RECT 34.456 65.536 51.378 65.625 ;
        RECT 34.41 65.582 51.332 65.671 ;
        RECT 34.364 65.628 51.286 65.717 ;
        RECT 34.318 65.674 51.24 65.763 ;
        RECT 34.272 65.72 51.194 65.809 ;
        RECT 34.226 65.766 51.148 65.855 ;
        RECT 34.18 65.812 51.102 65.901 ;
        RECT 34.134 65.858 51.056 65.947 ;
        RECT 34.088 65.904 51.01 65.993 ;
        RECT 34.042 65.95 50.964 66.039 ;
        RECT 33.996 65.996 50.918 66.085 ;
        RECT 33.95 66.042 50.872 66.131 ;
        RECT 33.904 66.088 50.826 66.177 ;
        RECT 33.858 66.134 50.78 66.223 ;
        RECT 33.812 66.18 50.734 66.269 ;
        RECT 33.766 66.226 50.688 66.315 ;
        RECT 33.72 66.272 50.642 66.361 ;
        RECT 33.674 66.318 50.596 66.407 ;
        RECT 33.628 66.364 50.55 66.453 ;
        RECT 33.582 66.41 50.504 66.499 ;
        RECT 33.536 66.456 50.458 66.545 ;
        RECT 33.49 66.502 50.412 66.591 ;
        RECT 33.444 66.548 50.366 66.637 ;
        RECT 33.398 66.594 50.32 66.683 ;
        RECT 33.352 66.64 50.274 66.729 ;
        RECT 33.306 66.686 50.228 66.775 ;
        RECT 33.26 66.732 50.182 66.821 ;
        RECT 33.214 66.778 50.136 66.867 ;
        RECT 33.168 66.824 50.09 66.913 ;
        RECT 33.122 66.87 50.044 66.959 ;
        RECT 33.076 66.916 49.998 67.005 ;
        RECT 33.03 66.962 49.952 67.051 ;
        RECT 32.984 67.008 49.906 67.097 ;
        RECT 32.938 67.054 49.86 67.143 ;
        RECT 32.892 67.1 49.814 67.189 ;
        RECT 32.846 67.146 49.768 67.235 ;
        RECT 32.8 67.192 49.722 67.281 ;
        RECT 32.754 67.238 49.676 67.327 ;
        RECT 32.708 67.284 49.63 67.373 ;
        RECT 32.662 67.33 49.584 67.419 ;
        RECT 32.616 67.376 49.538 67.465 ;
        RECT 32.57 67.422 49.492 67.511 ;
        RECT 32.524 67.468 49.446 67.557 ;
        RECT 32.478 67.514 49.4 67.603 ;
        RECT 32.432 67.56 49.354 67.649 ;
        RECT 32.386 67.606 49.308 67.695 ;
        RECT 32.34 67.652 49.262 67.741 ;
        RECT 32.294 67.698 49.216 67.787 ;
        RECT 32.248 67.744 49.17 67.833 ;
        RECT 32.202 67.79 49.124 67.879 ;
        RECT 32.156 67.836 49.078 67.925 ;
        RECT 32.11 67.882 49.032 67.971 ;
        RECT 32.064 67.928 48.986 68.017 ;
        RECT 32.018 67.974 48.94 68.063 ;
        RECT 31.972 68.02 48.894 68.109 ;
        RECT 31.926 68.066 48.848 68.155 ;
        RECT 31.88 68.112 48.802 68.201 ;
        RECT 31.834 68.158 48.756 68.247 ;
        RECT 31.788 68.204 48.71 68.293 ;
        RECT 31.742 68.25 48.664 68.339 ;
        RECT 31.696 68.296 48.618 68.385 ;
        RECT 31.65 68.342 48.572 68.431 ;
        RECT 31.604 68.388 48.526 68.477 ;
        RECT 31.558 68.434 48.48 68.523 ;
        RECT 31.512 68.48 48.434 68.569 ;
        RECT 31.466 68.526 48.388 68.615 ;
        RECT 31.42 68.572 48.342 68.661 ;
        RECT 31.374 68.618 48.296 68.707 ;
        RECT 31.328 68.664 48.25 68.753 ;
        RECT 31.282 68.71 48.204 68.799 ;
        RECT 31.236 68.756 48.158 68.845 ;
        RECT 31.19 68.802 48.112 68.891 ;
        RECT 31.144 68.848 48.066 68.937 ;
        RECT 31.098 68.894 48.02 68.983 ;
        RECT 31.052 68.94 47.974 69.029 ;
        RECT 31.006 68.986 47.928 69.075 ;
        RECT 30.96 69.032 47.882 69.121 ;
        RECT 30.914 69.078 47.836 69.167 ;
        RECT 30.868 69.124 47.79 69.213 ;
        RECT 30.822 69.17 47.744 69.259 ;
        RECT 30.776 69.216 47.698 69.305 ;
        RECT 30.73 69.262 47.652 69.351 ;
        RECT 30.684 69.308 47.606 69.397 ;
        RECT 30.638 69.354 47.56 69.443 ;
        RECT 30.592 69.4 47.514 69.489 ;
        RECT 30.546 69.446 47.468 69.535 ;
        RECT 30.5 69.492 47.422 69.581 ;
        RECT 30.5 69.492 47.376 69.627 ;
        RECT 30.5 69.492 47.33 69.673 ;
        RECT 30.5 69.492 47.284 69.719 ;
        RECT 30.5 69.492 47.238 69.765 ;
        RECT 30.5 69.492 47.192 69.811 ;
        RECT 30.5 69.492 47.146 69.857 ;
        RECT 30.5 69.492 47.1 69.903 ;
        RECT 30.5 69.492 47.054 69.949 ;
        RECT 30.5 69.492 47.008 69.995 ;
        RECT 30.5 69.492 46.962 70.041 ;
        RECT 30.5 69.492 46.916 70.087 ;
        RECT 30.5 69.492 46.87 70.133 ;
        RECT 30.5 69.492 46.824 70.179 ;
        RECT 30.5 69.492 46.778 70.225 ;
        RECT 30.5 69.492 46.732 70.271 ;
        RECT 30.5 69.492 46.686 70.317 ;
        RECT 30.5 69.492 46.64 70.363 ;
        RECT 30.5 69.492 46.594 70.409 ;
        RECT 30.5 69.492 46.548 70.455 ;
        RECT 30.5 69.492 46.502 70.501 ;
        RECT 30.5 69.492 46.456 70.547 ;
        RECT 30.5 69.492 46.41 70.593 ;
        RECT 30.5 69.492 46.364 70.639 ;
        RECT 30.5 69.492 46.318 70.685 ;
        RECT 30.5 69.492 46.272 70.731 ;
        RECT 30.5 69.492 46.226 70.777 ;
        RECT 30.5 69.492 46.18 70.823 ;
        RECT 30.5 69.492 46.134 70.869 ;
        RECT 30.5 69.492 46.088 70.915 ;
        RECT 30.5 69.492 46.042 70.961 ;
        RECT 30.5 69.492 45.996 71.007 ;
        RECT 30.5 69.492 45.95 71.053 ;
        RECT 30.5 69.492 45.904 71.099 ;
        RECT 30.5 69.492 45.858 71.145 ;
        RECT 30.5 69.492 45.812 71.191 ;
        RECT 30.5 69.492 45.766 71.237 ;
        RECT 30.5 69.492 45.72 71.283 ;
        RECT 30.5 69.492 45.674 71.329 ;
        RECT 30.5 69.492 45.628 71.375 ;
        RECT 30.5 69.492 45.582 71.421 ;
        RECT 30.5 69.492 45.536 71.467 ;
        RECT 30.5 69.492 45.49 71.513 ;
        RECT 30.5 69.492 45.444 71.559 ;
        RECT 30.5 69.492 45.398 71.605 ;
        RECT 30.5 69.492 45.352 71.651 ;
        RECT 30.5 69.492 45.306 71.697 ;
        RECT 30.5 69.492 45.26 71.743 ;
        RECT 30.5 69.492 45.214 71.789 ;
        RECT 30.5 69.492 45.168 71.835 ;
        RECT 30.5 69.492 45.122 71.881 ;
        RECT 30.5 69.492 45.076 71.927 ;
        RECT 30.5 69.492 45.03 71.973 ;
        RECT 30.5 69.492 44.984 72.019 ;
        RECT 30.5 69.492 44.938 72.065 ;
        RECT 30.5 69.492 44.892 72.111 ;
        RECT 30.5 69.492 44.846 72.157 ;
        RECT 30.5 69.492 44.8 72.203 ;
        RECT 30.5 69.492 44.754 72.249 ;
        RECT 30.5 69.492 44.708 72.295 ;
        RECT 30.5 69.492 44.662 72.341 ;
        RECT 30.5 69.492 44.616 72.387 ;
        RECT 30.5 69.492 44.57 72.433 ;
        RECT 30.5 69.492 44.524 72.479 ;
        RECT 30.5 69.492 44.478 72.525 ;
        RECT 30.5 69.492 44.432 72.571 ;
        RECT 30.5 69.492 44.386 72.617 ;
        RECT 30.5 69.492 44.34 72.663 ;
        RECT 30.5 69.492 44.294 72.709 ;
        RECT 30.5 69.492 44.248 72.755 ;
        RECT 30.5 69.492 44.202 72.801 ;
        RECT 30.5 69.492 44.156 72.847 ;
        RECT 30.5 69.492 44.11 72.893 ;
        RECT 30.5 69.492 44.064 72.939 ;
        RECT 30.5 69.492 44.018 72.985 ;
        RECT 30.5 69.492 43.972 73.031 ;
        RECT 30.5 69.492 43.926 73.077 ;
        RECT 30.5 69.492 43.88 73.123 ;
        RECT 30.5 69.492 43.834 73.169 ;
        RECT 30.5 69.492 43.788 73.215 ;
        RECT 30.5 69.492 43.742 73.261 ;
        RECT 30.5 69.492 43.696 73.307 ;
        RECT 30.5 69.492 43.65 73.353 ;
        RECT 30.5 69.492 43.604 73.399 ;
        RECT 30.5 69.492 43.558 73.445 ;
        RECT 30.5 69.492 43.512 73.491 ;
        RECT 30.5 69.492 43.466 73.537 ;
        RECT 30.5 69.492 43.42 73.583 ;
        RECT 30.5 69.492 43.374 73.629 ;
        RECT 30.5 69.492 43.328 73.675 ;
        RECT 30.5 69.492 43.282 73.721 ;
        RECT 30.5 69.492 43.236 73.767 ;
        RECT 30.5 69.492 43.19 73.813 ;
        RECT 30.5 69.492 43.144 73.859 ;
        RECT 30.5 69.492 43.098 73.905 ;
        RECT 30.5 69.492 43.052 73.951 ;
        RECT 30.5 69.492 43.006 73.997 ;
        RECT 30.5 69.492 42.96 74.043 ;
        RECT 30.5 69.492 42.914 74.089 ;
        RECT 30.5 69.492 42.868 74.135 ;
        RECT 30.5 69.492 42.822 74.181 ;
        RECT 30.5 69.492 42.776 74.227 ;
        RECT 30.5 69.492 42.73 74.273 ;
        RECT 30.5 69.492 42.684 74.319 ;
        RECT 30.5 69.492 42.638 74.365 ;
        RECT 30.5 69.492 42.592 74.411 ;
        RECT 30.5 69.492 42.546 74.457 ;
        RECT 30.5 69.492 42.5 110 ;
        RECT 76.265 44 110 56 ;
        RECT 59.312 60.93 76.265 60.978 ;
        RECT 59.358 60.884 76.311 60.942 ;
        RECT 76.24 44.012 76.265 60.978 ;
        RECT 59.404 60.838 76.357 60.896 ;
        RECT 76.194 44.048 76.24 61.013 ;
        RECT 59.266 60.976 76.194 61.059 ;
        RECT 59.45 60.792 76.403 60.85 ;
        RECT 76.148 44.094 76.194 61.059 ;
        RECT 59.22 61.022 76.148 61.105 ;
        RECT 59.496 60.746 76.449 60.804 ;
        RECT 76.102 44.14 76.148 61.105 ;
        RECT 59.174 61.068 76.102 61.151 ;
        RECT 59.542 60.7 76.495 60.758 ;
        RECT 76.056 44.186 76.102 61.151 ;
        RECT 59.128 61.114 76.056 61.197 ;
        RECT 59.588 60.654 76.541 60.712 ;
        RECT 76.01 44.232 76.056 61.197 ;
        RECT 59.082 61.16 76.01 61.243 ;
        RECT 59.634 60.608 76.587 60.666 ;
        RECT 75.964 44.278 76.01 61.243 ;
        RECT 59.036 61.206 75.964 61.289 ;
        RECT 59.68 60.562 76.633 60.62 ;
        RECT 75.918 44.324 75.964 61.289 ;
        RECT 58.99 61.252 75.918 61.335 ;
        RECT 59.726 60.516 76.679 60.574 ;
        RECT 75.872 44.37 75.918 61.335 ;
        RECT 58.944 61.298 75.872 61.381 ;
        RECT 59.772 60.47 76.725 60.528 ;
        RECT 75.826 44.416 75.872 61.381 ;
        RECT 58.898 61.344 75.826 61.427 ;
        RECT 59.818 60.424 76.771 60.482 ;
        RECT 75.78 44.462 75.826 61.427 ;
        RECT 58.852 61.39 75.78 61.473 ;
        RECT 59.864 60.378 76.817 60.436 ;
        RECT 75.734 44.508 75.78 61.473 ;
        RECT 58.806 61.436 75.734 61.519 ;
        RECT 59.91 60.332 76.863 60.39 ;
        RECT 75.688 44.554 75.734 61.519 ;
        RECT 58.76 61.482 75.688 61.565 ;
        RECT 59.956 60.286 76.909 60.344 ;
        RECT 75.642 44.6 75.688 61.565 ;
      LAYER MET4 ;
        RECT 70.814 69.423 79.278 69.485 ;
        RECT 77.852 62.385 110 63.5 ;
        RECT 79.232 61.005 79.278 69.485 ;
        RECT 70.768 69.469 79.232 69.531 ;
        RECT 77.898 62.339 110 63.5 ;
        RECT 79.186 61.051 79.232 69.531 ;
        RECT 70.722 69.515 79.186 69.577 ;
        RECT 77.944 62.293 110 63.5 ;
        RECT 79.14 61.097 79.186 69.577 ;
        RECT 70.676 69.561 79.14 69.623 ;
        RECT 77.99 62.247 110 63.5 ;
        RECT 79.094 61.143 79.14 69.623 ;
        RECT 70.63 69.607 79.094 69.669 ;
        RECT 78.036 62.201 110 63.5 ;
        RECT 79.048 61.189 79.094 69.669 ;
        RECT 70.584 69.653 79.048 69.715 ;
        RECT 78.082 62.155 110 63.5 ;
        RECT 79.002 61.235 79.048 69.715 ;
        RECT 70.538 69.699 79.002 69.761 ;
        RECT 78.128 62.109 110 63.5 ;
        RECT 78.956 61.281 79.002 69.761 ;
        RECT 70.492 69.745 78.956 69.807 ;
        RECT 78.174 62.063 110 63.5 ;
        RECT 78.91 61.327 78.956 69.807 ;
        RECT 70.446 69.791 78.91 69.853 ;
        RECT 78.22 62.017 110 63.5 ;
        RECT 78.864 61.373 78.91 69.853 ;
        RECT 70.4 69.837 78.864 69.899 ;
        RECT 78.266 61.971 110 63.5 ;
        RECT 78.818 61.419 78.864 69.899 ;
        RECT 70.354 69.883 78.818 69.945 ;
        RECT 78.312 61.925 110 63.5 ;
        RECT 78.772 61.465 78.818 69.945 ;
        RECT 70.308 69.929 78.772 69.991 ;
        RECT 78.358 61.879 110 63.5 ;
        RECT 78.726 61.511 78.772 69.991 ;
        RECT 70.262 69.975 78.726 70.037 ;
        RECT 78.404 61.833 110 63.5 ;
        RECT 78.68 61.557 78.726 70.037 ;
        RECT 70.216 70.021 78.68 70.083 ;
        RECT 78.45 61.787 110 63.5 ;
        RECT 78.634 61.603 78.68 70.083 ;
        RECT 70.17 70.067 78.634 70.129 ;
        RECT 78.496 61.741 110 63.5 ;
        RECT 78.588 61.649 78.634 70.129 ;
        RECT 70.124 70.113 78.588 70.175 ;
        RECT 78.542 61.695 110 63.5 ;
        RECT 70.078 70.159 78.542 70.221 ;
        RECT 70.032 70.205 78.496 70.267 ;
        RECT 69.986 70.251 78.45 70.313 ;
        RECT 69.94 70.297 78.404 70.359 ;
        RECT 69.894 70.343 78.358 70.405 ;
        RECT 69.848 70.389 78.312 70.451 ;
        RECT 69.802 70.435 78.266 70.497 ;
        RECT 69.756 70.481 78.22 70.543 ;
        RECT 69.71 70.527 78.174 70.589 ;
        RECT 69.664 70.573 78.128 70.635 ;
        RECT 69.618 70.619 78.082 70.681 ;
        RECT 69.572 70.665 78.036 70.727 ;
        RECT 69.526 70.711 77.99 70.773 ;
        RECT 69.48 70.757 77.944 70.819 ;
        RECT 69.434 70.803 77.898 70.865 ;
        RECT 69.388 70.849 77.852 70.911 ;
        RECT 69.342 70.895 77.806 70.957 ;
        RECT 69.296 70.941 77.76 71.003 ;
        RECT 69.25 70.987 77.714 71.049 ;
        RECT 69.204 71.033 77.668 71.095 ;
        RECT 69.158 71.079 77.622 71.141 ;
        RECT 69.112 71.125 77.576 71.187 ;
        RECT 69.066 71.171 77.53 71.233 ;
        RECT 69.02 71.217 77.484 71.279 ;
        RECT 68.974 71.263 77.438 71.325 ;
        RECT 68.928 71.309 77.392 71.371 ;
        RECT 68.882 71.355 77.346 71.417 ;
        RECT 68.836 71.401 77.3 71.463 ;
        RECT 68.79 71.447 77.254 71.509 ;
        RECT 68.744 71.493 77.208 71.555 ;
        RECT 68.698 71.539 77.162 71.601 ;
        RECT 68.652 71.585 77.116 71.647 ;
        RECT 68.606 71.631 77.07 71.693 ;
        RECT 68.56 71.677 77.024 71.739 ;
        RECT 68.514 71.723 76.978 71.785 ;
        RECT 68.468 71.769 76.932 71.831 ;
        RECT 68.422 71.815 76.886 71.877 ;
        RECT 68.376 71.861 76.84 71.923 ;
        RECT 68.33 71.907 76.794 71.969 ;
        RECT 68.284 71.953 76.748 72.015 ;
        RECT 68.238 71.999 76.702 72.061 ;
        RECT 68.192 72.045 76.656 72.107 ;
        RECT 68.146 72.091 76.61 72.153 ;
        RECT 68.1 72.137 76.564 72.199 ;
        RECT 68.054 72.183 76.518 72.245 ;
        RECT 68.008 72.229 76.472 72.291 ;
        RECT 67.962 72.275 76.426 72.337 ;
        RECT 67.916 72.321 76.38 72.383 ;
        RECT 67.87 72.367 76.334 72.429 ;
        RECT 67.824 72.413 76.288 72.475 ;
        RECT 67.778 72.459 76.242 72.521 ;
        RECT 67.732 72.505 76.196 72.567 ;
        RECT 67.686 72.551 76.15 72.613 ;
        RECT 67.64 72.597 76.104 72.659 ;
        RECT 67.594 72.643 76.058 72.705 ;
        RECT 67.548 72.689 76.012 72.751 ;
        RECT 67.502 72.735 75.966 72.797 ;
        RECT 67.456 72.781 75.92 72.843 ;
        RECT 67.41 72.827 75.874 72.889 ;
        RECT 67.364 72.873 75.828 72.935 ;
        RECT 67.318 72.919 75.782 72.981 ;
        RECT 67.272 72.965 75.736 73.027 ;
        RECT 67.226 73.011 75.69 73.073 ;
        RECT 67.18 73.057 75.644 73.119 ;
        RECT 67.134 73.103 75.598 73.165 ;
        RECT 67.088 73.149 75.552 73.211 ;
        RECT 67.042 73.195 75.506 73.257 ;
        RECT 66.996 73.241 75.46 73.303 ;
        RECT 66.95 73.287 75.414 73.349 ;
        RECT 66.904 73.333 75.368 73.395 ;
        RECT 66.858 73.379 75.322 73.441 ;
        RECT 66.812 73.425 75.276 73.487 ;
        RECT 66.766 73.471 75.23 73.533 ;
        RECT 66.72 73.517 75.184 73.579 ;
        RECT 66.674 73.563 75.138 73.625 ;
        RECT 66.628 73.609 75.092 73.671 ;
        RECT 66.582 73.655 75.046 73.717 ;
        RECT 66.536 73.701 75 73.763 ;
        RECT 66.49 73.747 74.954 73.809 ;
        RECT 66.444 73.793 74.908 73.855 ;
        RECT 66.398 73.839 74.862 73.901 ;
        RECT 66.352 73.885 74.816 73.947 ;
        RECT 66.306 73.931 74.77 73.993 ;
        RECT 66.26 73.977 74.724 74.039 ;
        RECT 66.214 74.023 74.678 74.085 ;
        RECT 66.168 74.069 74.632 74.131 ;
        RECT 66.122 74.115 74.586 74.177 ;
        RECT 66.076 74.161 74.54 74.223 ;
        RECT 66.03 74.207 74.494 74.269 ;
        RECT 65.984 74.253 74.448 74.315 ;
        RECT 65.938 74.299 74.402 74.361 ;
        RECT 65.892 74.345 74.356 74.407 ;
        RECT 65.846 74.391 74.31 74.453 ;
        RECT 65.8 74.437 74.264 74.499 ;
        RECT 65.754 74.483 74.218 74.545 ;
        RECT 65.708 74.529 74.172 74.591 ;
        RECT 65.662 74.575 74.126 74.637 ;
        RECT 65.616 74.621 74.08 74.683 ;
        RECT 65.57 74.667 74.034 74.729 ;
        RECT 65.524 74.713 73.988 74.775 ;
        RECT 65.478 74.759 73.942 74.821 ;
        RECT 65.432 74.805 73.896 74.867 ;
        RECT 65.386 74.851 73.85 74.913 ;
        RECT 65.34 74.897 73.804 74.959 ;
        RECT 65.294 74.943 73.758 75.005 ;
        RECT 65.248 74.989 73.712 75.051 ;
        RECT 65.202 75.035 73.666 75.097 ;
        RECT 65.156 75.081 73.62 75.143 ;
        RECT 65.11 75.127 73.574 75.189 ;
        RECT 65.064 75.173 73.528 75.235 ;
        RECT 65.018 75.219 73.482 75.281 ;
        RECT 64.972 75.265 73.436 75.327 ;
        RECT 64.926 75.311 73.39 75.373 ;
        RECT 64.88 75.357 73.344 75.419 ;
        RECT 64.834 75.403 73.298 75.465 ;
        RECT 64.788 75.449 73.252 75.511 ;
        RECT 64.742 75.495 73.206 75.557 ;
        RECT 64.696 75.541 73.16 75.603 ;
        RECT 64.65 75.587 73.114 75.649 ;
        RECT 64.604 75.633 73.068 75.695 ;
        RECT 64.558 75.679 73.022 75.741 ;
        RECT 64.512 75.725 72.976 75.787 ;
        RECT 64.466 75.771 72.93 75.833 ;
        RECT 64.42 75.817 72.884 75.879 ;
        RECT 64.374 75.863 72.838 75.925 ;
        RECT 64.328 75.909 72.792 75.971 ;
        RECT 64.282 75.955 72.746 76.017 ;
        RECT 64.236 76.001 72.7 76.063 ;
        RECT 64.19 76.047 72.654 76.109 ;
        RECT 64.144 76.093 72.608 76.155 ;
        RECT 64.098 76.139 72.562 76.201 ;
        RECT 64.052 76.185 72.516 76.247 ;
        RECT 64.006 76.231 72.47 76.293 ;
        RECT 63.96 76.277 72.424 76.339 ;
        RECT 63.914 76.323 72.378 76.385 ;
        RECT 63.868 76.369 72.332 76.431 ;
        RECT 63.822 76.415 72.286 76.477 ;
        RECT 63.776 76.461 72.24 76.523 ;
        RECT 63.73 76.507 72.194 76.569 ;
        RECT 63.684 76.553 72.148 76.615 ;
        RECT 63.638 76.599 72.102 76.661 ;
        RECT 63.592 76.645 72.056 76.707 ;
        RECT 63.546 76.691 72.01 76.753 ;
        RECT 63.5 76.737 71.964 76.799 ;
        RECT 63.48 76.77 71.918 76.845 ;
        RECT 63.434 76.803 71.872 76.891 ;
        RECT 63.388 76.849 71.826 76.937 ;
        RECT 63.342 76.895 71.78 76.983 ;
        RECT 63.296 76.941 71.734 77.029 ;
        RECT 63.25 76.987 71.688 77.075 ;
        RECT 63.204 77.033 71.642 77.121 ;
        RECT 63.158 77.079 71.596 77.167 ;
        RECT 63.112 77.125 71.55 77.213 ;
        RECT 63.066 77.171 71.504 77.259 ;
        RECT 63.02 77.217 71.458 77.305 ;
        RECT 62.974 77.263 71.412 77.351 ;
        RECT 62.928 77.309 71.366 77.397 ;
        RECT 62.882 77.355 71.32 77.443 ;
        RECT 62.836 77.401 71.274 77.489 ;
        RECT 62.79 77.447 71.228 77.535 ;
        RECT 62.744 77.493 71.182 77.581 ;
        RECT 62.698 77.539 71.136 77.627 ;
        RECT 62.652 77.585 71.09 77.673 ;
        RECT 62.606 77.631 71.044 77.719 ;
        RECT 62.56 77.677 70.998 77.765 ;
        RECT 62.514 77.723 70.952 77.811 ;
        RECT 62.468 77.769 70.906 77.857 ;
        RECT 62.422 77.815 70.86 77.903 ;
        RECT 62.376 77.861 70.814 77.949 ;
        RECT 62.33 77.907 70.768 77.995 ;
        RECT 62.284 77.953 70.722 78.041 ;
        RECT 62.238 77.999 70.676 78.087 ;
        RECT 62.192 78.045 70.63 78.133 ;
        RECT 62.146 78.091 70.584 78.179 ;
        RECT 62.1 78.137 70.538 78.225 ;
        RECT 62.054 78.183 70.492 78.271 ;
        RECT 62.008 78.229 70.446 78.317 ;
        RECT 61.962 78.275 70.4 78.363 ;
        RECT 61.916 78.321 70.354 78.409 ;
        RECT 61.87 78.367 70.308 78.455 ;
        RECT 61.824 78.413 70.262 78.501 ;
        RECT 61.778 78.459 70.216 78.547 ;
        RECT 61.732 78.505 70.17 78.593 ;
        RECT 61.686 78.551 70.124 78.639 ;
        RECT 61.64 78.597 70.078 78.685 ;
        RECT 61.594 78.643 70.032 78.731 ;
        RECT 61.548 78.689 69.986 78.777 ;
        RECT 61.502 78.735 69.94 78.823 ;
        RECT 61.456 78.781 69.894 78.869 ;
        RECT 61.41 78.827 69.848 78.915 ;
        RECT 61.364 78.873 69.802 78.961 ;
        RECT 61.318 78.919 69.756 79.007 ;
        RECT 61.272 78.965 69.71 79.053 ;
        RECT 61.226 79.011 69.664 79.099 ;
        RECT 61.18 79.057 69.618 79.145 ;
        RECT 61.134 79.103 69.572 79.191 ;
        RECT 61.088 79.149 69.526 79.237 ;
        RECT 61.042 79.195 69.48 79.283 ;
        RECT 60.996 79.241 69.434 79.329 ;
        RECT 60.95 79.287 69.388 79.375 ;
        RECT 60.904 79.333 69.342 79.421 ;
        RECT 60.858 79.379 69.296 79.467 ;
        RECT 60.812 79.425 69.25 79.513 ;
        RECT 60.766 79.471 69.204 79.559 ;
        RECT 60.72 79.517 69.158 79.605 ;
        RECT 60.674 79.563 69.112 79.651 ;
        RECT 60.628 79.609 69.066 79.697 ;
        RECT 60.582 79.655 69.02 79.743 ;
        RECT 60.536 79.701 68.974 79.789 ;
        RECT 60.49 79.747 68.928 79.835 ;
        RECT 60.444 79.793 68.882 79.881 ;
        RECT 60.398 79.839 68.836 79.927 ;
        RECT 60.352 79.885 68.79 79.973 ;
        RECT 60.306 79.931 68.744 80.019 ;
        RECT 60.26 79.977 68.698 80.065 ;
        RECT 60.214 80.023 68.652 80.111 ;
        RECT 60.168 80.069 68.606 80.157 ;
        RECT 60.122 80.115 68.56 80.203 ;
        RECT 60.076 80.161 68.514 80.249 ;
        RECT 60.03 80.207 68.468 80.295 ;
        RECT 59.984 80.253 68.422 80.341 ;
        RECT 59.938 80.299 68.376 80.387 ;
        RECT 59.892 80.345 68.33 80.433 ;
        RECT 59.846 80.391 68.284 80.479 ;
        RECT 59.8 80.437 68.238 80.525 ;
        RECT 59.754 80.483 68.192 80.571 ;
        RECT 59.708 80.529 68.146 80.617 ;
        RECT 59.662 80.575 68.1 80.663 ;
        RECT 59.616 80.621 68.054 80.709 ;
        RECT 59.57 80.667 68.008 80.755 ;
        RECT 59.524 80.713 67.962 80.801 ;
        RECT 59.478 80.759 67.916 80.847 ;
        RECT 59.432 80.805 67.87 80.893 ;
        RECT 59.386 80.851 67.824 80.939 ;
        RECT 59.34 80.897 67.778 80.985 ;
        RECT 59.294 80.943 67.732 81.031 ;
        RECT 59.248 80.989 67.686 81.077 ;
        RECT 59.202 81.035 67.64 81.123 ;
        RECT 59.156 81.081 67.594 81.169 ;
        RECT 59.11 81.127 67.548 81.215 ;
        RECT 59.064 81.173 67.502 81.261 ;
        RECT 59.018 81.219 67.456 81.307 ;
        RECT 58.972 81.265 67.41 81.353 ;
        RECT 58.926 81.311 67.364 81.399 ;
        RECT 58.88 81.357 67.318 81.445 ;
        RECT 58.834 81.403 67.272 81.491 ;
        RECT 58.788 81.449 67.226 81.537 ;
        RECT 58.742 81.495 67.18 81.583 ;
        RECT 58.696 81.541 67.134 81.629 ;
        RECT 58.65 81.587 67.088 81.675 ;
        RECT 58.604 81.633 67.042 81.721 ;
        RECT 58.558 81.679 66.996 81.767 ;
        RECT 58.512 81.725 66.95 81.813 ;
        RECT 58.466 81.771 66.904 81.859 ;
        RECT 58.42 81.817 66.858 81.905 ;
        RECT 58.374 81.863 66.812 81.951 ;
        RECT 58.328 81.909 66.766 81.997 ;
        RECT 58.282 81.955 66.72 82.043 ;
        RECT 58.236 82.001 66.674 82.089 ;
        RECT 58.19 82.047 66.628 82.135 ;
        RECT 58.144 82.093 66.582 82.181 ;
        RECT 58.098 82.139 66.536 82.227 ;
        RECT 58.052 82.185 66.49 82.273 ;
        RECT 58.006 82.231 66.444 82.319 ;
        RECT 57.96 82.277 66.398 82.365 ;
        RECT 57.914 82.323 66.352 82.411 ;
        RECT 57.868 82.369 66.306 82.457 ;
        RECT 57.822 82.415 66.26 82.503 ;
        RECT 57.776 82.461 66.214 82.549 ;
        RECT 57.73 82.507 66.168 82.595 ;
        RECT 57.684 82.553 66.122 82.641 ;
        RECT 57.638 82.599 66.076 82.687 ;
        RECT 57.592 82.645 66.03 82.733 ;
        RECT 57.546 82.691 65.984 82.779 ;
        RECT 57.5 82.737 65.938 82.825 ;
        RECT 57.5 82.737 65.892 82.871 ;
        RECT 57.5 82.737 65.846 82.917 ;
        RECT 57.5 82.737 65.8 82.963 ;
        RECT 57.5 82.737 65.754 83.009 ;
        RECT 57.5 82.737 65.708 83.055 ;
        RECT 57.5 82.737 65.662 83.101 ;
        RECT 57.5 82.737 65.616 83.147 ;
        RECT 57.5 82.737 65.57 83.193 ;
        RECT 57.5 82.737 65.524 83.239 ;
        RECT 57.5 82.737 65.478 83.285 ;
        RECT 57.5 82.737 65.432 83.331 ;
        RECT 57.5 82.737 65.386 83.377 ;
        RECT 57.5 82.737 65.34 83.423 ;
        RECT 57.5 82.737 65.294 83.469 ;
        RECT 57.5 82.737 65.248 83.515 ;
        RECT 57.5 82.737 65.202 83.561 ;
        RECT 57.5 82.737 65.156 83.607 ;
        RECT 57.5 82.737 65.11 83.653 ;
        RECT 57.5 82.737 65.064 83.699 ;
        RECT 57.5 82.737 65.018 83.745 ;
        RECT 57.5 82.737 64.972 83.791 ;
        RECT 57.5 82.737 64.926 83.837 ;
        RECT 57.5 82.737 64.88 83.883 ;
        RECT 57.5 82.737 64.834 83.929 ;
        RECT 57.5 82.737 64.788 83.975 ;
        RECT 57.5 82.737 64.742 84.021 ;
        RECT 57.5 82.737 64.696 84.067 ;
        RECT 57.5 82.737 64.65 84.113 ;
        RECT 57.5 82.737 64.604 84.159 ;
        RECT 57.5 82.737 64.558 84.205 ;
        RECT 57.5 82.737 64.512 84.251 ;
        RECT 57.5 82.737 64.466 84.297 ;
        RECT 57.5 82.737 64.42 84.343 ;
        RECT 57.5 82.737 64.374 84.389 ;
        RECT 57.5 82.737 64.328 84.435 ;
        RECT 57.5 82.737 64.282 84.481 ;
        RECT 57.5 82.737 64.236 84.527 ;
        RECT 57.5 82.737 64.19 84.573 ;
        RECT 57.5 82.737 64.144 84.619 ;
        RECT 57.5 82.737 64.098 84.665 ;
        RECT 57.5 82.737 64.052 84.711 ;
        RECT 57.5 82.737 64.006 84.757 ;
        RECT 57.5 82.737 63.96 84.803 ;
        RECT 57.5 82.737 63.914 84.849 ;
        RECT 57.5 82.737 63.868 84.895 ;
        RECT 57.5 82.737 63.822 84.941 ;
        RECT 57.5 82.737 63.776 84.987 ;
        RECT 57.5 82.737 63.73 85.033 ;
        RECT 57.5 82.737 63.684 85.079 ;
        RECT 57.5 82.737 63.638 85.125 ;
        RECT 57.5 82.737 63.592 85.171 ;
        RECT 57.5 82.737 63.546 85.217 ;
        RECT 57.5 82.737 63.5 110 ;
        RECT 88.365 68.5 110 77 ;
        RECT 79.852 76.99 91.885 77.012 ;
        RECT 76.366 80.476 88.365 80.522 ;
        RECT 76.412 80.43 88.411 80.497 ;
        RECT 88.362 68.501 88.365 80.522 ;
        RECT 76.458 80.384 88.457 80.451 ;
        RECT 88.316 68.526 88.362 80.546 ;
        RECT 76.32 80.522 88.316 80.592 ;
        RECT 76.504 80.338 88.503 80.405 ;
        RECT 88.27 68.572 88.316 80.592 ;
        RECT 76.274 80.568 88.27 80.638 ;
        RECT 76.55 80.292 88.549 80.359 ;
        RECT 88.224 68.618 88.27 80.638 ;
        RECT 76.228 80.614 88.224 80.684 ;
        RECT 76.596 80.246 88.595 80.313 ;
        RECT 88.178 68.664 88.224 80.684 ;
        RECT 76.182 80.66 88.178 80.73 ;
        RECT 76.642 80.2 88.641 80.267 ;
        RECT 88.132 68.71 88.178 80.73 ;
        RECT 76.136 80.706 88.132 80.776 ;
        RECT 76.688 80.154 88.687 80.221 ;
        RECT 88.086 68.756 88.132 80.776 ;
        RECT 76.09 80.752 88.086 80.822 ;
        RECT 76.734 80.108 88.733 80.175 ;
        RECT 88.04 68.802 88.086 80.822 ;
        RECT 76.044 80.798 88.04 80.868 ;
        RECT 76.78 80.062 88.779 80.129 ;
        RECT 87.994 68.848 88.04 80.868 ;
        RECT 75.998 80.844 87.994 80.914 ;
        RECT 76.826 80.016 88.825 80.083 ;
        RECT 87.948 68.894 87.994 80.914 ;
        RECT 75.952 80.89 87.948 80.96 ;
        RECT 76.872 79.97 88.871 80.037 ;
        RECT 87.902 68.94 87.948 80.96 ;
        RECT 75.906 80.936 87.902 81.006 ;
        RECT 76.918 79.924 88.917 79.991 ;
        RECT 87.856 68.986 87.902 81.006 ;
        RECT 75.86 80.982 87.856 81.052 ;
        RECT 76.964 79.883 88.963 79.945 ;
        RECT 87.81 69.032 87.856 81.052 ;
        RECT 75.814 81.028 87.81 81.098 ;
        RECT 77 79.842 89.009 79.899 ;
        RECT 87.764 69.078 87.81 81.098 ;
        RECT 75.768 81.074 87.764 81.144 ;
        RECT 77.046 79.796 89.055 79.853 ;
        RECT 87.718 69.124 87.764 81.144 ;
        RECT 75.722 81.12 87.718 81.19 ;
        RECT 77.092 79.75 89.101 79.807 ;
        RECT 87.672 69.17 87.718 81.19 ;
        RECT 75.676 81.166 87.672 81.236 ;
        RECT 77.138 79.704 89.147 79.761 ;
        RECT 87.626 69.216 87.672 81.236 ;
        RECT 75.63 81.212 87.626 81.282 ;
        RECT 77.184 79.658 89.193 79.715 ;
        RECT 87.58 69.262 87.626 81.282 ;
        RECT 75.584 81.258 87.58 81.328 ;
        RECT 77.23 79.612 89.239 79.669 ;
        RECT 87.534 69.308 87.58 81.328 ;
        RECT 75.538 81.304 87.534 81.374 ;
        RECT 77.276 79.566 89.285 79.623 ;
        RECT 87.488 69.354 87.534 81.374 ;
        RECT 75.492 81.35 87.488 81.42 ;
        RECT 77.322 79.52 89.331 79.577 ;
        RECT 87.442 69.4 87.488 81.42 ;
        RECT 75.446 81.396 87.442 81.466 ;
        RECT 77.368 79.474 89.377 79.531 ;
        RECT 87.396 69.446 87.442 81.466 ;
        RECT 75.4 81.442 87.396 81.512 ;
        RECT 77.414 79.428 89.423 79.485 ;
        RECT 87.35 69.492 87.396 81.512 ;
        RECT 75.354 81.488 87.35 81.558 ;
        RECT 77.46 79.382 89.469 79.439 ;
        RECT 87.304 69.538 87.35 81.558 ;
        RECT 75.308 81.534 87.304 81.604 ;
        RECT 77.506 79.336 89.515 79.393 ;
        RECT 87.258 69.584 87.304 81.604 ;
        RECT 75.262 81.58 87.258 81.65 ;
        RECT 77.552 79.29 89.561 79.347 ;
        RECT 87.212 69.63 87.258 81.65 ;
        RECT 75.216 81.626 87.212 81.696 ;
        RECT 77.598 79.244 89.607 79.301 ;
        RECT 87.166 69.676 87.212 81.696 ;
        RECT 75.17 81.672 87.166 81.742 ;
        RECT 77.644 79.198 89.653 79.255 ;
        RECT 87.12 69.722 87.166 81.742 ;
        RECT 75.124 81.718 87.12 81.788 ;
        RECT 77.69 79.152 89.699 79.209 ;
        RECT 87.074 69.768 87.12 81.788 ;
        RECT 75.078 81.764 87.074 81.834 ;
        RECT 77.736 79.106 89.745 79.163 ;
        RECT 87.028 69.814 87.074 81.834 ;
        RECT 75.032 81.81 87.028 81.88 ;
        RECT 77.782 79.06 89.791 79.117 ;
        RECT 86.982 69.86 87.028 81.88 ;
        RECT 74.986 81.856 86.982 81.926 ;
        RECT 77.828 79.014 89.837 79.071 ;
        RECT 86.936 69.906 86.982 81.926 ;
        RECT 74.94 81.902 86.936 81.972 ;
        RECT 77.874 78.968 89.883 79.025 ;
        RECT 86.89 69.952 86.936 81.972 ;
        RECT 74.894 81.948 86.89 82.018 ;
        RECT 77.92 78.922 89.929 78.979 ;
        RECT 86.844 69.998 86.89 82.018 ;
        RECT 74.848 81.994 86.844 82.064 ;
        RECT 77.966 78.876 89.975 78.933 ;
        RECT 86.798 70.044 86.844 82.064 ;
        RECT 74.802 82.04 86.798 82.11 ;
        RECT 78.012 78.83 90.021 78.887 ;
        RECT 86.752 70.09 86.798 82.11 ;
        RECT 74.756 82.086 86.752 82.156 ;
        RECT 78.058 78.784 90.067 78.841 ;
        RECT 86.706 70.136 86.752 82.156 ;
        RECT 74.71 82.132 86.706 82.202 ;
        RECT 78.104 78.738 90.113 78.795 ;
        RECT 86.66 70.182 86.706 82.202 ;
        RECT 74.664 82.178 86.66 82.248 ;
        RECT 78.15 78.692 90.159 78.749 ;
        RECT 86.614 70.228 86.66 82.248 ;
        RECT 74.618 82.224 86.614 82.294 ;
        RECT 78.196 78.646 90.205 78.703 ;
        RECT 86.568 70.274 86.614 82.294 ;
        RECT 74.572 82.27 86.568 82.34 ;
        RECT 78.242 78.6 90.251 78.657 ;
        RECT 86.522 70.32 86.568 82.34 ;
        RECT 74.526 82.316 86.522 82.386 ;
        RECT 78.288 78.554 90.297 78.611 ;
        RECT 86.476 70.366 86.522 82.386 ;
        RECT 74.48 82.362 86.476 82.432 ;
        RECT 78.334 78.508 90.343 78.565 ;
        RECT 86.43 70.412 86.476 82.432 ;
        RECT 74.434 82.408 86.43 82.478 ;
        RECT 78.38 78.462 90.389 78.519 ;
        RECT 86.384 70.458 86.43 82.478 ;
        RECT 74.388 82.454 86.384 82.524 ;
        RECT 78.426 78.416 90.435 78.473 ;
        RECT 86.338 70.504 86.384 82.524 ;
        RECT 74.342 82.5 86.338 82.57 ;
        RECT 78.472 78.37 90.481 78.427 ;
        RECT 86.292 70.55 86.338 82.57 ;
        RECT 74.296 82.546 86.292 82.616 ;
        RECT 78.518 78.324 90.527 78.381 ;
        RECT 86.246 70.596 86.292 82.616 ;
        RECT 74.25 82.592 86.246 82.662 ;
        RECT 78.564 78.278 90.573 78.335 ;
        RECT 86.2 70.642 86.246 82.662 ;
        RECT 74.204 82.638 86.2 82.708 ;
        RECT 78.61 78.232 90.619 78.289 ;
        RECT 86.154 70.688 86.2 82.708 ;
        RECT 74.158 82.684 86.154 82.754 ;
        RECT 78.656 78.186 90.665 78.243 ;
        RECT 86.108 70.734 86.154 82.754 ;
        RECT 74.112 82.73 86.108 82.8 ;
        RECT 78.702 78.14 90.711 78.197 ;
        RECT 86.062 70.78 86.108 82.8 ;
        RECT 74.066 82.776 86.062 82.846 ;
        RECT 78.748 78.094 90.757 78.151 ;
        RECT 86.016 70.826 86.062 82.846 ;
        RECT 74.02 82.822 86.016 82.892 ;
        RECT 78.794 78.048 90.803 78.105 ;
        RECT 85.97 70.872 86.016 82.892 ;
        RECT 73.974 82.868 85.97 82.938 ;
        RECT 78.84 78.002 90.849 78.059 ;
        RECT 85.924 70.918 85.97 82.938 ;
        RECT 73.928 82.914 85.924 82.984 ;
        RECT 78.886 77.956 90.895 78.013 ;
        RECT 85.878 70.964 85.924 82.984 ;
        RECT 73.882 82.96 85.878 83.03 ;
        RECT 78.932 77.91 90.941 77.967 ;
        RECT 85.832 71.01 85.878 83.03 ;
        RECT 73.836 83.006 85.832 83.076 ;
        RECT 78.978 77.864 90.987 77.921 ;
        RECT 85.786 71.056 85.832 83.076 ;
        RECT 73.79 83.052 85.786 83.122 ;
        RECT 79.024 77.818 91.033 77.875 ;
        RECT 85.74 71.102 85.786 83.122 ;
        RECT 73.744 83.098 85.74 83.168 ;
        RECT 79.07 77.772 91.079 77.829 ;
        RECT 85.694 71.148 85.74 83.168 ;
        RECT 73.698 83.144 85.694 83.214 ;
        RECT 79.116 77.726 91.125 77.783 ;
        RECT 85.648 71.194 85.694 83.214 ;
        RECT 73.652 83.19 85.648 83.26 ;
        RECT 79.162 77.68 91.171 77.737 ;
        RECT 85.602 71.24 85.648 83.26 ;
        RECT 73.606 83.236 85.602 83.306 ;
        RECT 79.208 77.634 91.217 77.691 ;
        RECT 85.556 71.286 85.602 83.306 ;
        RECT 73.56 83.282 85.556 83.352 ;
        RECT 79.254 77.588 91.263 77.645 ;
        RECT 85.51 71.332 85.556 83.352 ;
        RECT 73.514 83.328 85.51 83.398 ;
        RECT 79.3 77.542 91.309 77.599 ;
        RECT 85.464 71.378 85.51 83.398 ;
        RECT 73.468 83.374 85.464 83.444 ;
        RECT 79.346 77.496 91.355 77.553 ;
        RECT 85.418 71.424 85.464 83.444 ;
        RECT 73.422 83.42 85.418 83.49 ;
        RECT 79.392 77.45 91.401 77.507 ;
        RECT 85.372 71.47 85.418 83.49 ;
        RECT 73.376 83.466 85.372 83.536 ;
        RECT 79.438 77.404 91.447 77.461 ;
        RECT 85.326 71.516 85.372 83.536 ;
        RECT 73.33 83.512 85.326 83.582 ;
        RECT 79.484 77.358 91.493 77.415 ;
        RECT 85.28 71.562 85.326 83.582 ;
        RECT 73.284 83.558 85.28 83.628 ;
        RECT 79.53 77.312 91.539 77.369 ;
        RECT 85.234 71.608 85.28 83.628 ;
        RECT 73.238 83.604 85.234 83.674 ;
        RECT 79.576 77.266 91.585 77.323 ;
        RECT 85.188 71.654 85.234 83.674 ;
        RECT 73.192 83.65 85.188 83.72 ;
        RECT 79.622 77.22 91.631 77.277 ;
        RECT 85.142 71.7 85.188 83.72 ;
        RECT 73.146 83.696 85.142 83.766 ;
        RECT 79.668 77.174 91.677 77.231 ;
        RECT 85.096 71.746 85.142 83.766 ;
        RECT 73.1 83.742 85.096 83.812 ;
        RECT 79.714 77.128 91.723 77.185 ;
        RECT 85.05 71.792 85.096 83.812 ;
        RECT 73.054 83.788 85.05 83.858 ;
        RECT 79.76 77.082 91.769 77.139 ;
        RECT 85.004 71.838 85.05 83.858 ;
        RECT 73.008 83.834 85.004 83.904 ;
        RECT 79.806 77.036 91.815 77.093 ;
        RECT 84.958 71.884 85.004 83.904 ;
        RECT 72.962 83.88 84.958 83.95 ;
        RECT 79.852 76.99 91.861 77.047 ;
        RECT 84.912 71.93 84.958 83.95 ;
        RECT 72.916 83.926 84.912 83.996 ;
        RECT 79.898 76.944 110 77 ;
        RECT 84.866 71.976 84.912 83.996 ;
        RECT 72.87 83.972 84.866 84.042 ;
        RECT 79.944 76.898 110 77 ;
        RECT 84.82 72.022 84.866 84.042 ;
        RECT 72.824 84.018 84.82 84.088 ;
        RECT 79.99 76.852 110 77 ;
        RECT 84.774 72.068 84.82 84.088 ;
        RECT 72.778 84.064 84.774 84.134 ;
        RECT 80.036 76.806 110 77 ;
        RECT 84.728 72.114 84.774 84.134 ;
        RECT 72.732 84.11 84.728 84.18 ;
        RECT 80.082 76.76 110 77 ;
        RECT 84.682 72.16 84.728 84.18 ;
        RECT 72.686 84.156 84.682 84.226 ;
        RECT 80.128 76.714 110 77 ;
        RECT 84.636 72.206 84.682 84.226 ;
        RECT 72.64 84.202 84.636 84.272 ;
        RECT 80.174 76.668 110 77 ;
        RECT 84.59 72.252 84.636 84.272 ;
        RECT 72.594 84.248 84.59 84.318 ;
        RECT 80.22 76.622 110 77 ;
        RECT 84.544 72.298 84.59 84.318 ;
        RECT 72.548 84.294 84.544 84.364 ;
        RECT 80.266 76.576 110 77 ;
        RECT 84.498 72.344 84.544 84.364 ;
        RECT 72.502 84.34 84.498 84.41 ;
        RECT 80.312 76.53 110 77 ;
        RECT 84.452 72.39 84.498 84.41 ;
        RECT 72.456 84.386 84.452 84.456 ;
        RECT 80.358 76.484 110 77 ;
        RECT 84.406 72.436 84.452 84.456 ;
        RECT 72.41 84.432 84.406 84.502 ;
        RECT 80.404 76.438 110 77 ;
        RECT 84.36 72.482 84.406 84.502 ;
        RECT 72.364 84.478 84.36 84.548 ;
        RECT 80.45 76.392 110 77 ;
        RECT 84.314 72.528 84.36 84.548 ;
        RECT 72.318 84.524 84.314 84.594 ;
        RECT 80.496 76.346 110 77 ;
        RECT 84.268 72.574 84.314 84.594 ;
        RECT 72.272 84.57 84.268 84.64 ;
        RECT 80.542 76.3 110 77 ;
        RECT 84.222 72.62 84.268 84.64 ;
        RECT 72.226 84.616 84.222 84.686 ;
        RECT 80.588 76.254 110 77 ;
        RECT 84.176 72.666 84.222 84.686 ;
        RECT 72.18 84.662 84.176 84.732 ;
        RECT 80.634 76.208 110 77 ;
        RECT 84.13 72.712 84.176 84.732 ;
        RECT 72.134 84.708 84.13 84.778 ;
        RECT 80.68 76.162 110 77 ;
        RECT 84.084 72.758 84.13 84.778 ;
        RECT 72.088 84.754 84.084 84.824 ;
        RECT 80.726 76.116 110 77 ;
        RECT 84.038 72.804 84.084 84.824 ;
        RECT 72.042 84.8 84.038 84.87 ;
        RECT 80.772 76.07 110 77 ;
        RECT 83.992 72.85 84.038 84.87 ;
        RECT 71.996 84.846 83.992 84.916 ;
        RECT 80.818 76.024 110 77 ;
        RECT 83.946 72.896 83.992 84.916 ;
        RECT 71.95 84.892 83.946 84.962 ;
        RECT 80.864 75.978 110 77 ;
        RECT 83.9 72.942 83.946 84.962 ;
        RECT 71.904 84.938 83.9 85.008 ;
        RECT 80.91 75.932 110 77 ;
        RECT 83.854 72.988 83.9 85.008 ;
        RECT 71.858 84.984 83.854 85.054 ;
        RECT 80.956 75.886 110 77 ;
        RECT 83.808 73.034 83.854 85.054 ;
        RECT 71.812 85.03 83.808 85.1 ;
        RECT 81.002 75.84 110 77 ;
        RECT 83.762 73.08 83.808 85.1 ;
        RECT 71.766 85.076 83.762 85.146 ;
        RECT 81.048 75.794 110 77 ;
        RECT 83.716 73.126 83.762 85.146 ;
        RECT 71.72 85.122 83.716 85.192 ;
        RECT 81.094 75.748 110 77 ;
        RECT 83.67 73.172 83.716 85.192 ;
        RECT 71.674 85.168 83.67 85.238 ;
        RECT 81.14 75.702 110 77 ;
        RECT 83.624 73.218 83.67 85.238 ;
        RECT 71.628 85.214 83.624 85.284 ;
        RECT 81.186 75.656 110 77 ;
        RECT 83.578 73.264 83.624 85.284 ;
        RECT 71.582 85.26 83.578 85.33 ;
        RECT 81.232 75.61 110 77 ;
        RECT 83.532 73.31 83.578 85.33 ;
        RECT 71.536 85.306 83.532 85.376 ;
        RECT 81.278 75.564 110 77 ;
        RECT 83.486 73.356 83.532 85.376 ;
        RECT 71.49 85.352 83.486 85.422 ;
        RECT 81.324 75.518 110 77 ;
        RECT 83.44 73.402 83.486 85.422 ;
        RECT 71.444 85.398 83.44 85.468 ;
        RECT 81.37 75.472 110 77 ;
        RECT 83.394 73.448 83.44 85.468 ;
        RECT 71.398 85.444 83.394 85.514 ;
        RECT 81.416 75.426 110 77 ;
        RECT 83.348 73.494 83.394 85.514 ;
        RECT 71.352 85.49 83.348 85.56 ;
        RECT 81.462 75.38 110 77 ;
        RECT 83.302 73.54 83.348 85.56 ;
        RECT 71.306 85.536 83.302 85.606 ;
        RECT 81.508 75.334 110 77 ;
        RECT 83.256 73.586 83.302 85.606 ;
        RECT 71.26 85.582 83.256 85.652 ;
        RECT 81.554 75.288 110 77 ;
        RECT 83.21 73.632 83.256 85.652 ;
        RECT 71.214 85.628 83.21 85.698 ;
        RECT 81.6 75.242 110 77 ;
        RECT 83.164 73.678 83.21 85.698 ;
        RECT 71.168 85.674 83.164 85.744 ;
        RECT 81.646 75.196 110 77 ;
        RECT 83.118 73.724 83.164 85.744 ;
        RECT 71.122 85.72 83.118 85.79 ;
        RECT 81.692 75.15 110 77 ;
        RECT 83.072 73.77 83.118 85.79 ;
        RECT 71.076 85.766 83.072 85.836 ;
        RECT 81.738 75.104 110 77 ;
        RECT 83.026 73.816 83.072 85.836 ;
        RECT 71.03 85.812 83.026 85.882 ;
        RECT 81.784 75.058 110 77 ;
        RECT 82.98 73.862 83.026 85.882 ;
        RECT 70.984 85.858 82.98 85.928 ;
        RECT 81.83 75.012 110 77 ;
        RECT 82.934 73.908 82.98 85.928 ;
        RECT 70.938 85.904 82.934 85.974 ;
        RECT 81.876 74.966 110 77 ;
        RECT 82.888 73.954 82.934 85.974 ;
        RECT 70.892 85.95 82.888 86.02 ;
        RECT 81.922 74.92 110 77 ;
        RECT 82.842 74 82.888 86.02 ;
        RECT 70.846 85.996 82.842 86.066 ;
        RECT 81.968 74.874 110 77 ;
        RECT 82.796 74.046 82.842 86.066 ;
        RECT 70.8 86.042 82.796 86.112 ;
        RECT 82.014 74.828 110 77 ;
        RECT 82.75 74.092 82.796 86.112 ;
        RECT 70.754 86.088 82.75 86.158 ;
        RECT 82.06 74.782 110 77 ;
        RECT 82.704 74.138 82.75 86.158 ;
        RECT 70.708 86.134 82.704 86.204 ;
        RECT 82.106 74.736 110 77 ;
        RECT 82.658 74.184 82.704 86.204 ;
        RECT 70.662 86.18 82.658 86.25 ;
        RECT 82.152 74.69 110 77 ;
        RECT 82.612 74.23 82.658 86.25 ;
        RECT 70.616 86.226 82.612 86.296 ;
        RECT 82.198 74.644 110 77 ;
        RECT 82.566 74.276 82.612 86.296 ;
        RECT 70.57 86.272 82.566 86.342 ;
        RECT 82.244 74.598 110 77 ;
        RECT 82.52 74.322 82.566 86.342 ;
        RECT 70.524 86.318 82.52 86.388 ;
        RECT 82.29 74.552 110 77 ;
        RECT 82.474 74.368 82.52 86.388 ;
        RECT 70.478 86.364 82.474 86.434 ;
        RECT 82.336 74.506 110 77 ;
        RECT 82.428 74.414 82.474 86.434 ;
        RECT 70.432 86.41 82.428 86.48 ;
        RECT 82.382 74.46 110 77 ;
        RECT 70.386 86.456 82.382 86.526 ;
        RECT 70.34 86.502 82.336 86.572 ;
        RECT 70.294 86.548 82.29 86.618 ;
        RECT 70.248 86.594 82.244 86.664 ;
        RECT 70.202 86.64 82.198 86.71 ;
        RECT 70.156 86.686 82.152 86.756 ;
        RECT 70.11 86.732 82.106 86.802 ;
        RECT 70.064 86.778 82.06 86.848 ;
        RECT 70.018 86.824 82.014 86.894 ;
        RECT 69.972 86.87 81.968 86.94 ;
        RECT 69.926 86.916 81.922 86.986 ;
        RECT 69.88 86.962 81.876 87.032 ;
        RECT 69.834 87.008 81.83 87.078 ;
        RECT 69.788 87.054 81.784 87.124 ;
        RECT 69.742 87.1 81.738 87.17 ;
        RECT 69.696 87.146 81.692 87.216 ;
        RECT 69.65 87.192 81.646 87.262 ;
        RECT 69.604 87.238 81.6 87.308 ;
        RECT 69.558 87.284 81.554 87.354 ;
        RECT 69.512 87.33 81.508 87.4 ;
        RECT 69.466 87.376 81.462 87.446 ;
        RECT 69.42 87.422 81.416 87.492 ;
        RECT 69.374 87.468 81.37 87.538 ;
        RECT 69.328 87.514 81.324 87.584 ;
        RECT 69.282 87.56 81.278 87.63 ;
        RECT 69.236 87.606 81.232 87.676 ;
        RECT 69.19 87.652 81.186 87.722 ;
        RECT 69.144 87.698 81.14 87.768 ;
        RECT 69.098 87.744 81.094 87.814 ;
        RECT 69.052 87.79 81.048 87.86 ;
        RECT 69.006 87.836 81.002 87.906 ;
        RECT 68.96 87.882 80.956 87.952 ;
        RECT 68.914 87.928 80.91 87.998 ;
        RECT 68.868 87.974 80.864 88.044 ;
        RECT 68.822 88.02 80.818 88.09 ;
        RECT 68.776 88.066 80.772 88.136 ;
        RECT 68.73 88.112 80.726 88.182 ;
        RECT 68.684 88.158 80.68 88.228 ;
        RECT 68.638 88.204 80.634 88.274 ;
        RECT 68.592 88.25 80.588 88.32 ;
        RECT 68.546 88.296 80.542 88.366 ;
        RECT 68.5 88.342 80.496 88.412 ;
        RECT 68.5 88.342 80.45 88.458 ;
        RECT 68.5 88.342 80.404 88.504 ;
        RECT 68.5 88.342 80.358 88.55 ;
        RECT 68.5 88.342 80.312 88.596 ;
        RECT 68.5 88.342 80.266 88.642 ;
        RECT 68.5 88.342 80.22 88.688 ;
        RECT 68.5 88.342 80.174 88.734 ;
        RECT 68.5 88.342 80.128 88.78 ;
        RECT 68.5 88.342 80.082 88.826 ;
        RECT 68.5 88.342 80.036 88.872 ;
        RECT 68.5 88.342 79.99 88.918 ;
        RECT 68.5 88.342 79.944 88.964 ;
        RECT 68.5 88.342 79.898 89.01 ;
        RECT 68.5 88.342 79.852 89.056 ;
        RECT 68.5 88.342 79.806 89.102 ;
        RECT 68.5 88.342 79.76 89.148 ;
        RECT 68.5 88.342 79.714 89.194 ;
        RECT 68.5 88.342 79.668 89.24 ;
        RECT 68.5 88.342 79.622 89.286 ;
        RECT 68.5 88.342 79.576 89.332 ;
        RECT 68.5 88.342 79.53 89.378 ;
        RECT 68.5 88.342 79.484 89.424 ;
        RECT 68.5 88.342 79.438 89.47 ;
        RECT 68.5 88.342 79.392 89.516 ;
        RECT 68.5 88.342 79.346 89.562 ;
        RECT 68.5 88.342 79.3 89.608 ;
        RECT 68.5 88.342 79.254 89.654 ;
        RECT 68.5 88.342 79.208 89.7 ;
        RECT 68.5 88.342 79.162 89.746 ;
        RECT 68.5 88.342 79.116 89.792 ;
        RECT 68.5 88.342 79.07 89.838 ;
        RECT 68.5 88.342 79.024 89.884 ;
        RECT 68.5 88.342 78.978 89.93 ;
        RECT 68.5 88.342 78.932 89.976 ;
        RECT 68.5 88.342 78.886 90.022 ;
        RECT 68.5 88.342 78.84 90.068 ;
        RECT 68.5 88.342 78.794 90.114 ;
        RECT 68.5 88.342 78.748 90.16 ;
        RECT 68.5 88.342 78.702 90.206 ;
        RECT 68.5 88.342 78.656 90.252 ;
        RECT 68.5 88.342 78.61 90.298 ;
        RECT 68.5 88.342 78.564 90.344 ;
        RECT 68.5 88.342 78.518 90.39 ;
        RECT 68.5 88.342 78.472 90.436 ;
        RECT 68.5 88.342 78.426 90.482 ;
        RECT 68.5 88.342 78.38 90.528 ;
        RECT 68.5 88.342 78.334 90.574 ;
        RECT 68.5 88.342 78.288 90.62 ;
        RECT 68.5 88.342 78.242 90.666 ;
        RECT 68.5 88.342 78.196 90.712 ;
        RECT 68.5 88.342 78.15 90.758 ;
        RECT 68.5 88.342 78.104 90.804 ;
        RECT 68.5 88.342 78.058 90.85 ;
        RECT 68.5 88.342 78.012 90.896 ;
        RECT 68.5 88.342 77.966 90.942 ;
        RECT 68.5 88.342 77.92 90.988 ;
        RECT 68.5 88.342 77.874 91.034 ;
        RECT 68.5 88.342 77.828 91.08 ;
        RECT 68.5 88.342 77.782 91.126 ;
        RECT 68.5 88.342 77.736 91.172 ;
        RECT 68.5 88.342 77.69 91.218 ;
        RECT 68.5 88.342 77.644 91.264 ;
        RECT 68.5 88.342 77.598 91.31 ;
        RECT 68.5 88.342 77.552 91.356 ;
        RECT 68.5 88.342 77.506 91.402 ;
        RECT 68.5 88.342 77.46 91.448 ;
        RECT 68.5 88.342 77.414 91.494 ;
        RECT 68.5 88.342 77.368 91.54 ;
        RECT 68.5 88.342 77.322 91.586 ;
        RECT 68.5 88.342 77.276 91.632 ;
        RECT 68.5 88.342 77.23 91.678 ;
        RECT 68.5 88.342 77.184 91.724 ;
        RECT 68.5 88.342 77.138 91.77 ;
        RECT 68.5 88.342 77.092 91.816 ;
        RECT 68.5 88.342 77.046 91.862 ;
        RECT 68.5 88.342 77 110 ;
        RECT 75.642 44.6 75.688 61.57 ;
        RECT 58.714 61.528 75.642 61.616 ;
        RECT 60.002 60.24 76.955 60.303 ;
        RECT 75.596 44.646 75.642 61.616 ;
        RECT 58.668 61.574 75.596 61.662 ;
        RECT 60.048 60.194 77.001 60.257 ;
        RECT 75.55 44.692 75.596 61.662 ;
        RECT 58.622 61.62 75.55 61.708 ;
        RECT 60.094 60.148 77.047 60.211 ;
        RECT 75.504 44.738 75.55 61.708 ;
        RECT 58.576 61.666 75.504 61.754 ;
        RECT 60.14 60.102 77.093 60.165 ;
        RECT 75.458 44.784 75.504 61.754 ;
        RECT 58.53 61.712 75.458 61.8 ;
        RECT 60.186 60.056 77.139 60.119 ;
        RECT 75.412 44.83 75.458 61.8 ;
        RECT 58.484 61.758 75.412 61.846 ;
        RECT 60.232 60.01 77.185 60.073 ;
        RECT 75.366 44.876 75.412 61.846 ;
        RECT 58.438 61.804 75.366 61.892 ;
        RECT 60.278 59.964 77.231 60.027 ;
        RECT 75.32 44.922 75.366 61.892 ;
        RECT 58.392 61.85 75.32 61.938 ;
        RECT 60.324 59.918 77.277 59.981 ;
        RECT 75.274 44.968 75.32 61.938 ;
        RECT 58.346 61.896 75.274 61.984 ;
        RECT 60.37 59.872 77.323 59.935 ;
        RECT 75.228 45.014 75.274 61.984 ;
        RECT 58.3 61.942 75.228 62.03 ;
        RECT 60.416 59.826 77.369 59.889 ;
        RECT 75.182 45.06 75.228 62.03 ;
        RECT 58.254 61.988 75.182 62.076 ;
        RECT 60.462 59.78 77.415 59.843 ;
        RECT 75.136 45.106 75.182 62.076 ;
        RECT 58.208 62.034 75.136 62.122 ;
        RECT 60.508 59.734 77.461 59.797 ;
        RECT 75.09 45.152 75.136 62.122 ;
        RECT 58.162 62.08 75.09 62.168 ;
        RECT 60.554 59.688 77.507 59.751 ;
        RECT 75.044 45.198 75.09 62.168 ;
        RECT 58.116 62.126 75.044 62.214 ;
        RECT 60.6 59.642 77.553 59.705 ;
        RECT 74.998 45.244 75.044 62.214 ;
        RECT 58.07 62.172 74.998 62.26 ;
        RECT 60.646 59.596 77.599 59.659 ;
        RECT 74.952 45.29 74.998 62.26 ;
        RECT 58.024 62.218 74.952 62.306 ;
        RECT 60.692 59.55 77.645 59.613 ;
        RECT 74.906 45.336 74.952 62.306 ;
        RECT 57.978 62.264 74.906 62.352 ;
        RECT 60.738 59.504 77.691 59.567 ;
        RECT 74.86 45.382 74.906 62.352 ;
        RECT 57.932 62.31 74.86 62.398 ;
        RECT 60.784 59.458 77.737 59.521 ;
        RECT 74.814 45.428 74.86 62.398 ;
        RECT 57.886 62.356 74.814 62.444 ;
        RECT 60.83 59.412 77.783 59.475 ;
        RECT 74.768 45.474 74.814 62.444 ;
        RECT 57.84 62.402 74.768 62.49 ;
        RECT 60.876 59.366 77.829 59.429 ;
        RECT 74.722 45.52 74.768 62.49 ;
        RECT 57.794 62.448 74.722 62.536 ;
        RECT 60.922 59.32 77.875 59.383 ;
        RECT 74.676 45.566 74.722 62.536 ;
        RECT 57.748 62.494 74.676 62.582 ;
        RECT 60.968 59.274 77.921 59.337 ;
        RECT 74.63 45.612 74.676 62.582 ;
        RECT 57.702 62.54 74.63 62.628 ;
        RECT 61.014 59.228 77.967 59.291 ;
        RECT 74.584 45.658 74.63 62.628 ;
        RECT 57.656 62.586 74.584 62.674 ;
        RECT 61.06 59.182 78.013 59.245 ;
        RECT 74.538 45.704 74.584 62.674 ;
        RECT 57.61 62.632 74.538 62.72 ;
        RECT 61.106 59.136 78.059 59.199 ;
        RECT 74.492 45.75 74.538 62.72 ;
        RECT 57.564 62.678 74.492 62.766 ;
        RECT 61.152 59.09 78.105 59.153 ;
        RECT 74.446 45.796 74.492 62.766 ;
        RECT 57.518 62.724 74.446 62.812 ;
        RECT 61.198 59.044 78.151 59.107 ;
        RECT 74.4 45.842 74.446 62.812 ;
        RECT 57.472 62.77 74.4 62.858 ;
        RECT 61.244 58.998 78.197 59.061 ;
        RECT 74.354 45.888 74.4 62.858 ;
        RECT 57.426 62.816 74.354 62.904 ;
        RECT 61.29 58.952 78.243 59.015 ;
        RECT 74.308 45.934 74.354 62.904 ;
        RECT 57.38 62.862 74.308 62.95 ;
        RECT 61.336 58.906 78.289 58.969 ;
        RECT 74.262 45.98 74.308 62.95 ;
        RECT 57.334 62.908 74.262 62.996 ;
        RECT 61.382 58.86 78.335 58.923 ;
        RECT 74.216 46.026 74.262 62.996 ;
        RECT 57.288 62.954 74.216 63.042 ;
        RECT 61.428 58.814 78.381 58.877 ;
        RECT 74.17 46.072 74.216 63.042 ;
        RECT 57.242 63 74.17 63.088 ;
        RECT 61.474 58.768 78.427 58.831 ;
        RECT 74.124 46.118 74.17 63.088 ;
        RECT 57.196 63.046 74.124 63.134 ;
        RECT 61.52 58.722 78.473 58.785 ;
        RECT 74.078 46.164 74.124 63.134 ;
        RECT 57.15 63.092 74.078 63.18 ;
        RECT 61.566 58.676 78.519 58.739 ;
        RECT 74.032 46.21 74.078 63.18 ;
        RECT 57.104 63.138 74.032 63.226 ;
        RECT 61.612 58.63 78.565 58.693 ;
        RECT 73.986 46.256 74.032 63.226 ;
        RECT 57.058 63.184 73.986 63.272 ;
        RECT 61.658 58.584 78.611 58.647 ;
        RECT 73.94 46.302 73.986 63.272 ;
        RECT 57.012 63.23 73.94 63.318 ;
        RECT 61.704 58.538 78.657 58.601 ;
        RECT 73.894 46.348 73.94 63.318 ;
        RECT 56.966 63.276 73.894 63.364 ;
        RECT 61.75 58.492 78.703 58.555 ;
        RECT 73.848 46.394 73.894 63.364 ;
        RECT 56.92 63.322 73.848 63.41 ;
        RECT 61.796 58.446 78.749 58.509 ;
        RECT 73.802 46.44 73.848 63.41 ;
        RECT 56.874 63.368 73.802 63.456 ;
        RECT 61.842 58.4 78.795 58.463 ;
        RECT 73.756 46.486 73.802 63.456 ;
        RECT 56.828 63.414 73.756 63.502 ;
        RECT 61.888 58.354 78.841 58.417 ;
        RECT 73.71 46.532 73.756 63.502 ;
        RECT 56.782 63.46 73.71 63.548 ;
        RECT 61.934 58.308 78.887 58.371 ;
        RECT 73.664 46.578 73.71 63.548 ;
        RECT 56.736 63.506 73.664 63.594 ;
        RECT 61.98 58.262 78.933 58.325 ;
        RECT 73.618 46.624 73.664 63.594 ;
        RECT 56.69 63.552 73.618 63.64 ;
        RECT 62.026 58.216 78.979 58.279 ;
        RECT 73.572 46.67 73.618 63.64 ;
        RECT 56.644 63.598 73.572 63.686 ;
        RECT 62.072 58.17 79.025 58.233 ;
        RECT 73.526 46.716 73.572 63.686 ;
        RECT 56.598 63.644 73.526 63.732 ;
        RECT 62.118 58.124 79.071 58.187 ;
        RECT 73.48 46.762 73.526 63.732 ;
        RECT 56.552 63.69 73.48 63.778 ;
        RECT 62.164 58.078 79.117 58.141 ;
        RECT 73.434 46.808 73.48 63.778 ;
        RECT 56.506 63.736 73.434 63.824 ;
        RECT 62.21 58.032 79.163 58.095 ;
        RECT 73.388 46.854 73.434 63.824 ;
        RECT 56.46 63.782 73.388 63.87 ;
        RECT 62.256 57.986 79.209 58.049 ;
        RECT 73.342 46.9 73.388 63.87 ;
        RECT 56.414 63.828 73.342 63.916 ;
        RECT 62.302 57.94 79.255 58.003 ;
        RECT 73.296 46.946 73.342 63.916 ;
        RECT 56.368 63.874 73.296 63.962 ;
        RECT 62.348 57.894 79.301 57.957 ;
        RECT 73.25 46.992 73.296 63.962 ;
        RECT 56.322 63.92 73.25 64.008 ;
        RECT 62.394 57.848 79.347 57.911 ;
        RECT 73.204 47.038 73.25 64.008 ;
        RECT 56.276 63.966 73.204 64.054 ;
        RECT 62.44 57.802 79.393 57.865 ;
        RECT 73.158 47.084 73.204 64.054 ;
        RECT 56.23 64.012 73.158 64.1 ;
        RECT 62.486 57.756 79.439 57.819 ;
        RECT 73.112 47.13 73.158 64.1 ;
        RECT 56.184 64.058 73.112 64.146 ;
        RECT 62.532 57.71 79.485 57.773 ;
        RECT 73.066 47.176 73.112 64.146 ;
        RECT 56.138 64.104 73.066 64.192 ;
        RECT 62.578 57.664 79.531 57.727 ;
        RECT 73.02 47.222 73.066 64.192 ;
        RECT 56.092 64.15 73.02 64.238 ;
        RECT 62.624 57.618 79.577 57.681 ;
        RECT 72.974 47.268 73.02 64.238 ;
        RECT 56 64.242 72.974 64.284 ;
        RECT 56.046 64.196 72.974 64.284 ;
        RECT 62.67 57.572 79.623 57.635 ;
        RECT 72.928 47.314 72.974 64.284 ;
        RECT 55.96 64.285 72.928 64.33 ;
        RECT 62.716 57.526 79.669 57.589 ;
        RECT 72.882 47.36 72.928 64.33 ;
        RECT 55.914 64.328 72.882 64.376 ;
        RECT 62.762 57.48 79.715 57.543 ;
        RECT 72.836 47.406 72.882 64.376 ;
        RECT 55.868 64.374 72.836 64.422 ;
        RECT 62.808 57.434 79.761 57.497 ;
        RECT 72.79 47.452 72.836 64.422 ;
        RECT 55.822 64.42 72.79 64.468 ;
        RECT 62.854 57.388 79.807 57.451 ;
        RECT 72.744 47.498 72.79 64.468 ;
        RECT 55.776 64.466 72.744 64.514 ;
        RECT 62.9 57.342 79.853 57.405 ;
        RECT 72.698 47.544 72.744 64.514 ;
        RECT 55.73 64.512 72.698 64.56 ;
        RECT 62.946 57.296 79.899 57.359 ;
        RECT 72.652 47.59 72.698 64.56 ;
        RECT 55.684 64.558 72.652 64.606 ;
        RECT 62.992 57.25 79.945 57.313 ;
        RECT 72.606 47.636 72.652 64.606 ;
        RECT 55.638 64.604 72.606 64.652 ;
        RECT 63.038 57.204 79.991 57.267 ;
        RECT 72.56 47.682 72.606 64.652 ;
        RECT 55.592 64.65 72.56 64.698 ;
        RECT 63.084 57.158 80.037 57.221 ;
        RECT 72.514 47.728 72.56 64.698 ;
        RECT 55.546 64.696 72.514 64.744 ;
        RECT 63.13 57.112 80.083 57.175 ;
        RECT 72.468 47.774 72.514 64.744 ;
        RECT 55.5 64.742 72.468 64.79 ;
        RECT 63.176 57.066 80.129 57.129 ;
        RECT 72.422 47.82 72.468 64.79 ;
        RECT 55.454 64.788 72.422 64.836 ;
        RECT 63.222 57.02 80.175 57.083 ;
        RECT 72.376 47.866 72.422 64.836 ;
        RECT 55.408 64.834 72.376 64.882 ;
        RECT 63.268 56.974 80.221 57.037 ;
        RECT 72.33 47.912 72.376 64.882 ;
        RECT 55.362 64.88 72.33 64.928 ;
        RECT 63.314 56.928 80.267 56.991 ;
        RECT 72.284 47.958 72.33 64.928 ;
        RECT 55.316 64.926 72.284 64.974 ;
        RECT 63.36 56.882 80.313 56.945 ;
        RECT 72.238 48.004 72.284 64.974 ;
        RECT 55.27 64.972 72.238 65.02 ;
        RECT 63.406 56.836 80.359 56.899 ;
        RECT 72.192 48.05 72.238 65.02 ;
        RECT 55.224 65.018 72.192 65.066 ;
        RECT 63.452 56.79 80.405 56.853 ;
        RECT 72.146 48.096 72.192 65.066 ;
        RECT 55.178 65.064 72.146 65.112 ;
        RECT 63.498 56.744 80.451 56.807 ;
        RECT 72.1 48.142 72.146 65.112 ;
        RECT 55.132 65.11 72.1 65.158 ;
        RECT 63.544 56.698 80.497 56.761 ;
        RECT 72.054 48.188 72.1 65.158 ;
        RECT 55.086 65.156 72.054 65.204 ;
        RECT 63.59 56.652 80.543 56.715 ;
        RECT 72.008 48.234 72.054 65.204 ;
        RECT 55.04 65.202 72.008 65.25 ;
        RECT 63.636 56.606 80.589 56.669 ;
        RECT 71.962 48.28 72.008 65.25 ;
        RECT 54.994 65.248 71.962 65.296 ;
        RECT 63.682 56.56 80.635 56.623 ;
        RECT 71.916 48.326 71.962 65.296 ;
        RECT 54.948 65.294 71.916 65.342 ;
        RECT 63.728 56.514 80.681 56.577 ;
        RECT 71.87 48.372 71.916 65.342 ;
        RECT 54.902 65.34 71.87 65.388 ;
        RECT 63.774 56.468 80.727 56.531 ;
        RECT 71.824 48.418 71.87 65.388 ;
        RECT 54.856 65.386 71.824 65.434 ;
        RECT 63.82 56.422 80.773 56.485 ;
        RECT 71.778 48.464 71.824 65.434 ;
        RECT 54.81 65.432 71.778 65.48 ;
        RECT 63.866 56.376 80.819 56.439 ;
        RECT 71.732 48.51 71.778 65.48 ;
        RECT 54.764 65.478 71.732 65.526 ;
        RECT 63.912 56.33 80.865 56.393 ;
        RECT 71.686 48.556 71.732 65.526 ;
        RECT 54.718 65.524 71.686 65.572 ;
        RECT 63.958 56.284 80.911 56.347 ;
        RECT 71.64 48.602 71.686 65.572 ;
        RECT 54.672 65.57 71.64 65.618 ;
        RECT 64.004 56.238 80.957 56.301 ;
        RECT 71.594 48.648 71.64 65.618 ;
        RECT 54.626 65.616 71.594 65.664 ;
        RECT 64.05 56.192 81.003 56.255 ;
        RECT 71.548 48.694 71.594 65.664 ;
        RECT 54.58 65.662 71.548 65.71 ;
        RECT 64.096 56.146 81.049 56.209 ;
        RECT 71.502 48.74 71.548 65.71 ;
        RECT 54.534 65.708 71.502 65.756 ;
        RECT 64.142 56.1 81.095 56.163 ;
        RECT 71.456 48.786 71.502 65.756 ;
        RECT 54.488 65.754 71.456 65.802 ;
        RECT 64.188 56.054 81.141 56.117 ;
        RECT 71.41 48.832 71.456 65.802 ;
        RECT 54.442 65.8 71.41 65.848 ;
        RECT 64.234 56.008 81.187 56.071 ;
        RECT 71.364 48.878 71.41 65.848 ;
        RECT 54.396 65.846 71.364 65.894 ;
        RECT 64.28 55.962 81.233 56.024 ;
        RECT 71.318 48.924 71.364 65.894 ;
        RECT 54.35 65.892 71.318 65.94 ;
        RECT 64.326 55.916 110 56 ;
        RECT 71.272 48.97 71.318 65.94 ;
        RECT 54.304 65.938 71.272 65.986 ;
        RECT 64.372 55.87 110 56 ;
        RECT 71.226 49.016 71.272 65.986 ;
        RECT 54.258 65.984 71.226 66.032 ;
        RECT 64.418 55.824 110 56 ;
        RECT 71.18 49.062 71.226 66.032 ;
        RECT 54.212 66.03 71.18 66.078 ;
        RECT 64.464 55.778 110 56 ;
        RECT 71.134 49.108 71.18 66.078 ;
        RECT 54.166 66.076 71.134 66.124 ;
        RECT 64.51 55.732 110 56 ;
        RECT 71.088 49.154 71.134 66.124 ;
        RECT 54.12 66.122 71.088 66.17 ;
        RECT 64.556 55.686 110 56 ;
        RECT 71.042 49.2 71.088 66.17 ;
        RECT 54.074 66.168 71.042 66.216 ;
        RECT 64.602 55.64 110 56 ;
        RECT 70.996 49.246 71.042 66.216 ;
        RECT 54.028 66.214 70.996 66.262 ;
        RECT 64.648 55.594 110 56 ;
        RECT 70.95 49.292 70.996 66.262 ;
        RECT 53.982 66.26 70.95 66.308 ;
        RECT 64.694 55.548 110 56 ;
        RECT 70.904 49.338 70.95 66.308 ;
        RECT 53.936 66.306 70.904 66.354 ;
        RECT 64.74 55.502 110 56 ;
        RECT 70.858 49.384 70.904 66.354 ;
        RECT 53.89 66.352 70.858 66.4 ;
        RECT 64.786 55.456 110 56 ;
        RECT 70.812 49.43 70.858 66.4 ;
        RECT 53.844 66.398 70.812 66.446 ;
        RECT 64.832 55.41 110 56 ;
        RECT 70.766 49.476 70.812 66.446 ;
        RECT 53.798 66.444 70.766 66.492 ;
        RECT 64.878 55.364 110 56 ;
        RECT 70.72 49.522 70.766 66.492 ;
        RECT 53.752 66.49 70.72 66.538 ;
        RECT 64.924 55.318 110 56 ;
        RECT 70.674 49.568 70.72 66.538 ;
        RECT 53.706 66.536 70.674 66.584 ;
        RECT 64.97 55.272 110 56 ;
        RECT 70.628 49.614 70.674 66.584 ;
        RECT 53.66 66.582 70.628 66.63 ;
        RECT 65.016 55.226 110 56 ;
        RECT 70.582 49.66 70.628 66.63 ;
        RECT 53.614 66.628 70.582 66.676 ;
        RECT 65.062 55.18 110 56 ;
        RECT 70.536 49.706 70.582 66.676 ;
        RECT 53.568 66.674 70.536 66.722 ;
        RECT 65.108 55.134 110 56 ;
        RECT 70.49 49.752 70.536 66.722 ;
        RECT 53.522 66.72 70.49 66.768 ;
        RECT 65.154 55.088 110 56 ;
        RECT 70.444 49.798 70.49 66.768 ;
        RECT 53.476 66.766 70.444 66.814 ;
        RECT 65.2 55.042 110 56 ;
        RECT 70.398 49.844 70.444 66.814 ;
        RECT 53.43 66.812 70.398 66.86 ;
        RECT 65.246 54.996 110 56 ;
        RECT 70.352 49.89 70.398 66.86 ;
        RECT 53.384 66.858 70.352 66.906 ;
        RECT 65.292 54.95 110 56 ;
        RECT 70.306 49.936 70.352 66.906 ;
        RECT 53.338 66.904 70.306 66.952 ;
        RECT 65.338 54.904 110 56 ;
        RECT 70.26 49.982 70.306 66.952 ;
        RECT 53.292 66.95 70.26 66.998 ;
        RECT 65.384 54.858 110 56 ;
        RECT 70.214 50.028 70.26 66.998 ;
        RECT 53.246 66.996 70.214 67.044 ;
        RECT 65.43 54.812 110 56 ;
        RECT 70.168 50.074 70.214 67.044 ;
        RECT 53.2 67.042 70.168 67.09 ;
        RECT 65.476 54.766 110 56 ;
        RECT 70.122 50.12 70.168 67.09 ;
        RECT 53.154 67.088 70.122 67.136 ;
        RECT 65.522 54.72 110 56 ;
        RECT 70.076 50.166 70.122 67.136 ;
        RECT 53.108 67.134 70.076 67.182 ;
        RECT 65.568 54.674 110 56 ;
        RECT 70.03 50.212 70.076 67.182 ;
        RECT 53.062 67.18 70.03 67.228 ;
        RECT 65.614 54.628 110 56 ;
        RECT 69.984 50.258 70.03 67.228 ;
        RECT 53.016 67.226 69.984 67.274 ;
        RECT 65.66 54.582 110 56 ;
        RECT 69.938 50.304 69.984 67.274 ;
        RECT 52.97 67.272 69.938 67.32 ;
        RECT 65.706 54.536 110 56 ;
        RECT 69.892 50.35 69.938 67.32 ;
        RECT 52.924 67.318 69.892 67.366 ;
        RECT 65.752 54.49 110 56 ;
        RECT 69.846 50.396 69.892 67.366 ;
        RECT 52.878 67.364 69.846 67.412 ;
        RECT 65.798 54.444 110 56 ;
        RECT 69.8 50.442 69.846 67.412 ;
        RECT 52.832 67.41 69.8 67.458 ;
        RECT 65.844 54.398 110 56 ;
        RECT 69.754 50.488 69.8 67.458 ;
        RECT 52.786 67.456 69.754 67.504 ;
        RECT 65.89 54.352 110 56 ;
        RECT 69.708 50.534 69.754 67.504 ;
        RECT 52.74 67.502 69.708 67.55 ;
        RECT 65.936 54.306 110 56 ;
        RECT 69.662 50.58 69.708 67.55 ;
        RECT 52.694 67.548 69.662 67.596 ;
        RECT 65.982 54.26 110 56 ;
        RECT 69.616 50.626 69.662 67.596 ;
        RECT 52.648 67.594 69.616 67.642 ;
        RECT 66.028 54.214 110 56 ;
        RECT 69.57 50.672 69.616 67.642 ;
        RECT 52.602 67.64 69.57 67.688 ;
        RECT 66.074 54.168 110 56 ;
        RECT 69.524 50.718 69.57 67.688 ;
        RECT 52.556 67.686 69.524 67.734 ;
        RECT 66.12 54.122 110 56 ;
        RECT 69.478 50.764 69.524 67.734 ;
        RECT 52.51 67.732 69.478 67.78 ;
        RECT 66.166 54.076 110 56 ;
        RECT 69.432 50.81 69.478 67.78 ;
        RECT 52.464 67.778 69.432 67.826 ;
        RECT 66.212 54.03 110 56 ;
        RECT 69.386 50.856 69.432 67.826 ;
        RECT 52.418 67.824 69.386 67.872 ;
        RECT 66.258 53.984 110 56 ;
        RECT 69.34 50.902 69.386 67.872 ;
        RECT 52.372 67.87 69.34 67.918 ;
        RECT 66.304 53.938 110 56 ;
        RECT 69.294 50.948 69.34 67.918 ;
        RECT 52.326 67.916 69.294 67.964 ;
        RECT 66.35 53.892 110 56 ;
        RECT 69.248 50.994 69.294 67.964 ;
        RECT 52.28 67.962 69.248 68.01 ;
        RECT 66.396 53.846 110 56 ;
        RECT 69.202 51.04 69.248 68.01 ;
        RECT 52.234 68.008 69.202 68.056 ;
        RECT 66.442 53.8 110 56 ;
        RECT 69.156 51.086 69.202 68.056 ;
        RECT 52.188 68.054 69.156 68.102 ;
        RECT 66.488 53.754 110 56 ;
        RECT 69.11 51.132 69.156 68.102 ;
        RECT 52.142 68.1 69.11 68.148 ;
        RECT 66.534 53.708 110 56 ;
        RECT 69.064 51.178 69.11 68.148 ;
        RECT 52.096 68.146 69.064 68.194 ;
        RECT 66.58 53.662 110 56 ;
        RECT 69.018 51.224 69.064 68.194 ;
        RECT 52.05 68.192 69.018 68.24 ;
        RECT 66.626 53.616 110 56 ;
        RECT 68.972 51.27 69.018 68.24 ;
        RECT 52.004 68.238 68.972 68.286 ;
        RECT 66.672 53.57 110 56 ;
        RECT 68.926 51.316 68.972 68.286 ;
        RECT 51.958 68.284 68.926 68.332 ;
        RECT 66.718 53.524 110 56 ;
        RECT 68.88 51.362 68.926 68.332 ;
        RECT 51.912 68.33 68.88 68.378 ;
        RECT 66.764 53.478 110 56 ;
        RECT 68.834 51.408 68.88 68.378 ;
        RECT 51.866 68.376 68.834 68.424 ;
        RECT 66.81 53.432 110 56 ;
        RECT 68.788 51.454 68.834 68.424 ;
        RECT 51.82 68.422 68.788 68.47 ;
        RECT 66.856 53.386 110 56 ;
        RECT 68.742 51.5 68.788 68.47 ;
        RECT 51.774 68.468 68.742 68.516 ;
        RECT 66.902 53.34 110 56 ;
        RECT 68.696 51.546 68.742 68.516 ;
        RECT 51.728 68.514 68.696 68.562 ;
        RECT 66.948 53.294 110 56 ;
        RECT 68.65 51.592 68.696 68.562 ;
        RECT 51.682 68.56 68.65 68.608 ;
        RECT 66.994 53.248 110 56 ;
        RECT 68.604 51.638 68.65 68.608 ;
        RECT 51.636 68.606 68.604 68.654 ;
        RECT 67.04 53.202 110 56 ;
        RECT 68.558 51.684 68.604 68.654 ;
        RECT 51.59 68.652 68.558 68.7 ;
        RECT 67.086 53.156 110 56 ;
        RECT 68.512 51.73 68.558 68.7 ;
        RECT 51.544 68.698 68.512 68.746 ;
        RECT 67.132 53.11 110 56 ;
        RECT 68.466 51.776 68.512 68.746 ;
        RECT 51.498 68.744 68.466 68.792 ;
        RECT 67.178 53.064 110 56 ;
        RECT 68.42 51.822 68.466 68.792 ;
        RECT 51.452 68.79 68.42 68.838 ;
        RECT 67.224 53.018 110 56 ;
        RECT 68.374 51.868 68.42 68.838 ;
        RECT 51.406 68.836 68.374 68.884 ;
        RECT 67.27 52.972 110 56 ;
        RECT 68.328 51.914 68.374 68.884 ;
        RECT 51.36 68.882 68.328 68.93 ;
        RECT 67.316 52.926 110 56 ;
        RECT 68.282 51.96 68.328 68.93 ;
        RECT 51.314 68.928 68.282 68.976 ;
        RECT 67.362 52.88 110 56 ;
        RECT 68.236 52.006 68.282 68.976 ;
        RECT 51.268 68.974 68.236 69.022 ;
        RECT 67.408 52.834 110 56 ;
        RECT 68.19 52.052 68.236 69.022 ;
        RECT 51.222 69.02 68.19 69.068 ;
        RECT 67.454 52.788 110 56 ;
        RECT 68.144 52.098 68.19 69.068 ;
        RECT 51.176 69.066 68.144 69.114 ;
        RECT 67.5 52.742 110 56 ;
        RECT 68.098 52.144 68.144 69.114 ;
        RECT 51.13 69.112 68.098 69.16 ;
        RECT 67.546 52.696 110 56 ;
        RECT 68.052 52.19 68.098 69.16 ;
        RECT 51.084 69.158 68.052 69.206 ;
        RECT 67.592 52.65 110 56 ;
        RECT 68.006 52.236 68.052 69.206 ;
        RECT 51.038 69.204 68.006 69.252 ;
        RECT 67.638 52.604 110 56 ;
        RECT 67.96 52.282 68.006 69.252 ;
        RECT 50.992 69.25 67.96 69.298 ;
        RECT 67.684 52.558 110 56 ;
        RECT 67.914 52.328 67.96 69.298 ;
        RECT 50.946 69.296 67.914 69.344 ;
        RECT 67.73 52.512 110 56 ;
        RECT 67.868 52.374 67.914 69.344 ;
        RECT 50.9 69.342 67.868 69.39 ;
        RECT 67.776 52.466 110 56 ;
        RECT 67.822 52.42 67.868 69.39 ;
        RECT 50.854 69.388 67.822 69.436 ;
        RECT 50.808 69.434 67.776 69.482 ;
        RECT 50.762 69.48 67.73 69.528 ;
        RECT 50.716 69.526 67.684 69.574 ;
        RECT 50.67 69.572 67.638 69.62 ;
        RECT 50.624 69.618 67.592 69.666 ;
        RECT 50.578 69.664 67.546 69.712 ;
        RECT 50.532 69.71 67.5 69.758 ;
        RECT 50.486 69.756 67.454 69.804 ;
        RECT 50.44 69.802 67.408 69.85 ;
        RECT 50.394 69.848 67.362 69.896 ;
        RECT 50.348 69.894 67.316 69.942 ;
        RECT 50.302 69.94 67.27 69.988 ;
        RECT 50.256 69.986 67.224 70.034 ;
        RECT 50.21 70.032 67.178 70.08 ;
        RECT 50.164 70.078 67.132 70.126 ;
        RECT 50.118 70.124 67.086 70.172 ;
        RECT 50.072 70.17 67.04 70.218 ;
        RECT 50.026 70.216 66.994 70.264 ;
        RECT 49.98 70.262 66.948 70.31 ;
        RECT 49.934 70.308 66.902 70.356 ;
        RECT 49.888 70.354 66.856 70.402 ;
        RECT 49.842 70.4 66.81 70.448 ;
        RECT 49.796 70.446 66.764 70.494 ;
        RECT 49.75 70.492 66.718 70.54 ;
        RECT 49.704 70.538 66.672 70.586 ;
        RECT 49.658 70.584 66.626 70.632 ;
        RECT 49.612 70.63 66.58 70.678 ;
        RECT 49.566 70.676 66.534 70.724 ;
        RECT 49.52 70.722 66.488 70.77 ;
        RECT 49.474 70.768 66.442 70.816 ;
        RECT 49.428 70.814 66.396 70.862 ;
        RECT 49.382 70.86 66.35 70.908 ;
        RECT 49.336 70.906 66.304 70.954 ;
        RECT 49.29 70.952 66.258 71 ;
        RECT 49.244 70.998 66.212 71.046 ;
        RECT 49.198 71.044 66.166 71.092 ;
        RECT 49.152 71.09 66.12 71.138 ;
        RECT 49.106 71.136 66.074 71.184 ;
        RECT 49.06 71.182 66.028 71.23 ;
        RECT 49.014 71.228 65.982 71.276 ;
        RECT 48.968 71.274 65.936 71.322 ;
        RECT 48.922 71.32 65.89 71.368 ;
        RECT 48.876 71.366 65.844 71.414 ;
        RECT 48.83 71.412 65.798 71.46 ;
        RECT 48.784 71.458 65.752 71.506 ;
        RECT 48.738 71.504 65.706 71.552 ;
        RECT 48.692 71.55 65.66 71.598 ;
        RECT 48.646 71.596 65.614 71.644 ;
        RECT 48.6 71.642 65.568 71.69 ;
        RECT 48.554 71.688 65.522 71.736 ;
        RECT 48.508 71.734 65.476 71.782 ;
        RECT 48.462 71.78 65.43 71.828 ;
        RECT 48.416 71.826 65.384 71.874 ;
        RECT 48.37 71.872 65.338 71.92 ;
        RECT 48.324 71.918 65.292 71.966 ;
        RECT 48.278 71.964 65.246 72.012 ;
        RECT 48.232 72.01 65.2 72.058 ;
        RECT 48.186 72.056 65.154 72.104 ;
        RECT 48.14 72.102 65.108 72.15 ;
        RECT 48.094 72.148 65.062 72.196 ;
        RECT 48.048 72.194 65.016 72.242 ;
        RECT 48.002 72.24 64.97 72.288 ;
        RECT 47.956 72.286 64.924 72.334 ;
        RECT 47.91 72.332 64.878 72.38 ;
        RECT 47.864 72.378 64.832 72.426 ;
        RECT 47.818 72.424 64.786 72.472 ;
        RECT 47.772 72.47 64.74 72.518 ;
        RECT 47.726 72.516 64.694 72.564 ;
        RECT 47.68 72.562 64.648 72.61 ;
        RECT 47.634 72.608 64.602 72.656 ;
        RECT 47.588 72.654 64.556 72.702 ;
        RECT 47.542 72.7 64.51 72.748 ;
        RECT 47.496 72.746 64.464 72.794 ;
        RECT 47.45 72.792 64.418 72.84 ;
        RECT 47.404 72.838 64.372 72.886 ;
        RECT 47.358 72.884 64.326 72.932 ;
        RECT 47.312 72.93 64.28 72.978 ;
        RECT 47.266 72.976 64.234 73.024 ;
        RECT 47.22 73.022 64.188 73.07 ;
        RECT 47.174 73.068 64.142 73.116 ;
        RECT 47.128 73.114 64.096 73.162 ;
        RECT 47.082 73.16 64.05 73.208 ;
        RECT 47.036 73.206 64.004 73.254 ;
        RECT 46.99 73.252 63.958 73.3 ;
        RECT 46.944 73.298 63.912 73.346 ;
        RECT 46.898 73.344 63.866 73.392 ;
        RECT 46.852 73.39 63.82 73.438 ;
        RECT 46.806 73.436 63.774 73.484 ;
        RECT 46.76 73.482 63.728 73.53 ;
        RECT 46.714 73.528 63.682 73.576 ;
        RECT 46.668 73.574 63.636 73.622 ;
        RECT 46.622 73.62 63.59 73.668 ;
        RECT 46.576 73.666 63.544 73.714 ;
        RECT 46.53 73.712 63.498 73.76 ;
        RECT 46.484 73.758 63.452 73.806 ;
        RECT 46.438 73.804 63.406 73.852 ;
        RECT 46.392 73.85 63.36 73.898 ;
        RECT 46.346 73.896 63.314 73.944 ;
        RECT 46.3 73.942 63.268 73.99 ;
        RECT 46.254 73.988 63.222 74.036 ;
        RECT 46.208 74.034 63.176 74.082 ;
        RECT 46.162 74.08 63.13 74.128 ;
        RECT 46.116 74.126 63.084 74.174 ;
        RECT 46.07 74.172 63.038 74.22 ;
        RECT 46.024 74.218 62.992 74.266 ;
        RECT 45.978 74.264 62.946 74.312 ;
        RECT 45.932 74.31 62.9 74.358 ;
        RECT 45.886 74.356 62.854 74.404 ;
        RECT 45.84 74.402 62.808 74.45 ;
        RECT 45.794 74.448 62.762 74.496 ;
        RECT 45.748 74.494 62.716 74.542 ;
        RECT 45.702 74.54 62.67 74.588 ;
        RECT 45.656 74.586 62.624 74.634 ;
        RECT 45.61 74.632 62.578 74.68 ;
        RECT 45.564 74.678 62.532 74.726 ;
        RECT 45.518 74.724 62.486 74.772 ;
        RECT 45.472 74.77 62.44 74.818 ;
        RECT 45.426 74.816 62.394 74.864 ;
        RECT 45.38 74.862 62.348 74.91 ;
        RECT 45.334 74.908 62.302 74.956 ;
        RECT 45.288 74.954 62.256 75.002 ;
        RECT 45.242 75 62.21 75.048 ;
        RECT 45.196 75.046 62.164 75.094 ;
        RECT 45.15 75.092 62.118 75.14 ;
        RECT 45.104 75.138 62.072 75.186 ;
        RECT 45.058 75.184 62.026 75.232 ;
        RECT 45.012 75.23 61.98 75.278 ;
        RECT 44.966 75.276 61.934 75.324 ;
        RECT 44.92 75.322 61.888 75.37 ;
        RECT 44.874 75.368 61.842 75.416 ;
        RECT 44.828 75.414 61.796 75.462 ;
        RECT 44.782 75.46 61.75 75.508 ;
        RECT 44.736 75.506 61.704 75.554 ;
        RECT 44.69 75.552 61.658 75.6 ;
        RECT 44.644 75.598 61.612 75.646 ;
        RECT 44.598 75.644 61.566 75.692 ;
        RECT 44.552 75.69 61.52 75.738 ;
        RECT 44.506 75.736 61.474 75.784 ;
        RECT 44.46 75.782 61.428 75.83 ;
        RECT 44.414 75.828 61.382 75.876 ;
        RECT 44.368 75.874 61.336 75.922 ;
        RECT 44.322 75.92 61.29 75.968 ;
        RECT 44.276 75.966 61.244 76.014 ;
        RECT 44.23 76.012 61.198 76.06 ;
        RECT 44.184 76.058 61.152 76.106 ;
        RECT 44.138 76.104 61.106 76.152 ;
        RECT 44.092 76.15 61.06 76.198 ;
        RECT 44.046 76.196 61.014 76.244 ;
        RECT 44 76.242 60.968 76.29 ;
        RECT 44 76.242 60.922 76.336 ;
        RECT 44 76.242 60.876 76.382 ;
        RECT 44 76.242 60.83 76.428 ;
        RECT 44 76.242 60.784 76.474 ;
        RECT 44 76.242 60.738 76.52 ;
        RECT 44 76.242 60.692 76.566 ;
        RECT 44 76.242 60.646 76.612 ;
        RECT 44 76.242 60.6 76.658 ;
        RECT 44 76.242 60.554 76.704 ;
        RECT 44 76.242 60.508 76.75 ;
        RECT 44 76.242 60.462 76.796 ;
        RECT 44 76.242 60.416 76.842 ;
        RECT 44 76.242 60.37 76.888 ;
        RECT 44 76.242 60.324 76.934 ;
        RECT 44 76.242 60.278 76.98 ;
        RECT 44 76.242 60.232 77.026 ;
        RECT 44 76.242 60.186 77.072 ;
        RECT 44 76.242 60.14 77.118 ;
        RECT 44 76.242 60.094 77.164 ;
        RECT 44 76.242 60.048 77.21 ;
        RECT 44 76.242 60.002 77.256 ;
        RECT 44 76.242 59.956 77.302 ;
        RECT 44 76.242 59.91 77.348 ;
        RECT 44 76.242 59.864 77.394 ;
        RECT 44 76.242 59.818 77.44 ;
        RECT 44 76.242 59.772 77.486 ;
        RECT 44 76.242 59.726 77.532 ;
        RECT 44 76.242 59.68 77.578 ;
        RECT 44 76.242 59.634 77.624 ;
        RECT 44 76.242 59.588 77.67 ;
        RECT 44 76.242 59.542 77.716 ;
        RECT 44 76.242 59.496 77.762 ;
        RECT 44 76.242 59.45 77.808 ;
        RECT 44 76.242 59.404 77.854 ;
        RECT 44 76.242 59.358 77.9 ;
        RECT 44 76.242 59.312 77.946 ;
        RECT 44 76.242 59.266 77.992 ;
        RECT 44 76.242 59.22 78.038 ;
        RECT 44 76.242 59.174 78.084 ;
        RECT 44 76.242 59.128 78.13 ;
        RECT 44 76.242 59.082 78.176 ;
        RECT 44 76.242 59.036 78.222 ;
        RECT 44 76.242 58.99 78.268 ;
        RECT 44 76.242 58.944 78.314 ;
        RECT 44 76.242 58.898 78.36 ;
        RECT 44 76.242 58.852 78.406 ;
        RECT 44 76.242 58.806 78.452 ;
        RECT 44 76.242 58.76 78.498 ;
        RECT 44 76.242 58.714 78.544 ;
        RECT 44 76.242 58.668 78.59 ;
        RECT 44 76.242 58.622 78.636 ;
        RECT 44 76.242 58.576 78.682 ;
        RECT 44 76.242 58.53 78.728 ;
        RECT 44 76.242 58.484 78.774 ;
        RECT 44 76.242 58.438 78.82 ;
        RECT 44 76.242 58.392 78.866 ;
        RECT 44 76.242 58.346 78.912 ;
        RECT 44 76.242 58.3 78.958 ;
        RECT 44 76.242 58.254 79.004 ;
        RECT 44 76.242 58.208 79.05 ;
        RECT 44 76.242 58.162 79.096 ;
        RECT 44 76.242 58.116 79.142 ;
        RECT 44 76.242 58.07 79.188 ;
        RECT 44 76.242 58.024 79.234 ;
        RECT 44 76.242 57.978 79.28 ;
        RECT 44 76.242 57.932 79.326 ;
        RECT 44 76.242 57.886 79.372 ;
        RECT 44 76.242 57.84 79.418 ;
        RECT 44 76.242 57.794 79.464 ;
        RECT 44 76.242 57.748 79.51 ;
        RECT 44 76.242 57.702 79.556 ;
        RECT 44 76.242 57.656 79.602 ;
        RECT 44 76.242 57.61 79.648 ;
        RECT 44 76.242 57.564 79.694 ;
        RECT 44 76.242 57.518 79.74 ;
        RECT 44 76.242 57.472 79.786 ;
        RECT 44 76.242 57.426 79.832 ;
        RECT 44 76.242 57.38 79.878 ;
        RECT 44 76.242 57.334 79.924 ;
        RECT 44 76.242 57.288 79.97 ;
        RECT 44 76.242 57.242 80.016 ;
        RECT 44 76.242 57.196 80.062 ;
        RECT 44 76.242 57.15 80.108 ;
        RECT 44 76.242 57.104 80.154 ;
        RECT 44 76.242 57.058 80.2 ;
        RECT 44 76.242 57.012 80.246 ;
        RECT 44 76.242 56.966 80.292 ;
        RECT 44 76.242 56.92 80.338 ;
        RECT 44 76.242 56.874 80.384 ;
        RECT 44 76.242 56.828 80.43 ;
        RECT 44 76.242 56.782 80.476 ;
        RECT 44 76.242 56.736 80.522 ;
        RECT 44 76.242 56.69 80.568 ;
        RECT 44 76.242 56.644 80.614 ;
        RECT 44 76.242 56.598 80.66 ;
        RECT 44 76.242 56.552 80.706 ;
        RECT 44 76.242 56.506 80.752 ;
        RECT 44 76.242 56.46 80.798 ;
        RECT 44 76.242 56.414 80.844 ;
        RECT 44 76.242 56.368 80.89 ;
        RECT 44 76.242 56.322 80.936 ;
        RECT 44 76.242 56.276 80.982 ;
        RECT 44 76.242 56.23 81.028 ;
        RECT 44 76.242 56.184 81.074 ;
        RECT 44 76.242 56.138 81.12 ;
        RECT 44 76.242 56.092 81.166 ;
        RECT 44 76.242 56.046 81.212 ;
        RECT 44 76.242 56 110 ;
        RECT 82.76 57.5 110 63.5 ;
        RECT 76.748 63.489 85.24 63.521 ;
        RECT 74.31 65.927 82.76 65.996 ;
        RECT 74.356 65.881 82.806 65.957 ;
        RECT 82.728 57.516 82.76 65.996 ;
        RECT 74.264 65.973 82.728 66.035 ;
        RECT 74.402 65.835 82.852 65.911 ;
        RECT 82.682 57.555 82.728 66.035 ;
        RECT 74.218 66.019 82.682 66.081 ;
        RECT 74.448 65.789 82.898 65.865 ;
        RECT 82.636 57.601 82.682 66.081 ;
        RECT 74.172 66.065 82.636 66.127 ;
        RECT 74.494 65.743 82.944 65.819 ;
        RECT 82.59 57.647 82.636 66.127 ;
        RECT 74.126 66.111 82.59 66.173 ;
        RECT 74.54 65.697 82.99 65.773 ;
        RECT 82.544 57.693 82.59 66.173 ;
        RECT 74.08 66.157 82.544 66.219 ;
        RECT 74.586 65.651 83.036 65.727 ;
        RECT 82.498 57.739 82.544 66.219 ;
        RECT 74.034 66.203 82.498 66.265 ;
        RECT 74.632 65.605 83.082 65.681 ;
        RECT 82.452 57.785 82.498 66.265 ;
        RECT 73.988 66.249 82.452 66.311 ;
        RECT 74.678 65.559 83.128 65.635 ;
        RECT 82.406 57.831 82.452 66.311 ;
        RECT 73.942 66.295 82.406 66.357 ;
        RECT 74.724 65.513 83.174 65.589 ;
        RECT 82.36 57.877 82.406 66.357 ;
        RECT 73.896 66.341 82.36 66.403 ;
        RECT 74.77 65.467 83.22 65.543 ;
        RECT 82.314 57.923 82.36 66.403 ;
        RECT 73.85 66.387 82.314 66.449 ;
        RECT 74.816 65.421 83.266 65.497 ;
        RECT 82.268 57.969 82.314 66.449 ;
        RECT 73.804 66.433 82.268 66.495 ;
        RECT 74.862 65.375 83.312 65.451 ;
        RECT 82.222 58.015 82.268 66.495 ;
        RECT 73.758 66.479 82.222 66.541 ;
        RECT 74.908 65.329 83.358 65.405 ;
        RECT 82.176 58.061 82.222 66.541 ;
        RECT 73.712 66.525 82.176 66.587 ;
        RECT 74.954 65.283 83.404 65.359 ;
        RECT 82.13 58.107 82.176 66.587 ;
        RECT 73.666 66.571 82.13 66.633 ;
        RECT 75 65.237 83.45 65.313 ;
        RECT 82.084 58.153 82.13 66.633 ;
        RECT 73.62 66.617 82.084 66.679 ;
        RECT 75.046 65.191 83.496 65.267 ;
        RECT 82.038 58.199 82.084 66.679 ;
        RECT 73.574 66.663 82.038 66.725 ;
        RECT 75.092 65.145 83.542 65.221 ;
        RECT 81.992 58.245 82.038 66.725 ;
        RECT 73.528 66.709 81.992 66.771 ;
        RECT 75.138 65.099 83.588 65.175 ;
        RECT 81.946 58.291 81.992 66.771 ;
        RECT 73.482 66.755 81.946 66.817 ;
        RECT 75.184 65.053 83.634 65.129 ;
        RECT 81.9 58.337 81.946 66.817 ;
        RECT 73.436 66.801 81.9 66.863 ;
        RECT 75.23 65.007 83.68 65.083 ;
        RECT 81.854 58.383 81.9 66.863 ;
        RECT 73.39 66.847 81.854 66.909 ;
        RECT 75.276 64.961 83.726 65.037 ;
        RECT 81.808 58.429 81.854 66.909 ;
        RECT 73.344 66.893 81.808 66.955 ;
        RECT 75.322 64.915 83.772 64.991 ;
        RECT 81.762 58.475 81.808 66.955 ;
        RECT 73.298 66.939 81.762 67.001 ;
        RECT 75.368 64.869 83.818 64.945 ;
        RECT 81.716 58.521 81.762 67.001 ;
        RECT 73.252 66.985 81.716 67.047 ;
        RECT 75.414 64.823 83.864 64.899 ;
        RECT 81.67 58.567 81.716 67.047 ;
        RECT 73.206 67.031 81.67 67.093 ;
        RECT 75.46 64.777 83.91 64.853 ;
        RECT 81.624 58.613 81.67 67.093 ;
        RECT 73.16 67.077 81.624 67.139 ;
        RECT 75.506 64.731 83.956 64.807 ;
        RECT 81.578 58.659 81.624 67.139 ;
        RECT 73.114 67.123 81.578 67.185 ;
        RECT 75.552 64.685 84.002 64.761 ;
        RECT 81.532 58.705 81.578 67.185 ;
        RECT 73.068 67.169 81.532 67.231 ;
        RECT 75.598 64.639 84.048 64.715 ;
        RECT 81.486 58.751 81.532 67.231 ;
        RECT 73.022 67.215 81.486 67.277 ;
        RECT 75.644 64.593 84.094 64.669 ;
        RECT 81.44 58.797 81.486 67.277 ;
        RECT 72.976 67.261 81.44 67.323 ;
        RECT 75.69 64.547 84.14 64.623 ;
        RECT 81.394 58.843 81.44 67.323 ;
        RECT 72.93 67.307 81.394 67.369 ;
        RECT 75.736 64.501 84.186 64.577 ;
        RECT 81.348 58.889 81.394 67.369 ;
        RECT 72.884 67.353 81.348 67.415 ;
        RECT 75.782 64.455 84.232 64.531 ;
        RECT 81.302 58.935 81.348 67.415 ;
        RECT 72.838 67.399 81.302 67.461 ;
        RECT 75.828 64.409 84.278 64.485 ;
        RECT 81.256 58.981 81.302 67.461 ;
        RECT 72.792 67.445 81.256 67.507 ;
        RECT 75.874 64.363 84.324 64.439 ;
        RECT 81.21 59.027 81.256 67.507 ;
        RECT 72.746 67.491 81.21 67.553 ;
        RECT 75.92 64.317 84.37 64.393 ;
        RECT 81.164 59.073 81.21 67.553 ;
        RECT 72.7 67.537 81.164 67.599 ;
        RECT 75.966 64.271 84.416 64.347 ;
        RECT 81.118 59.119 81.164 67.599 ;
        RECT 72.654 67.583 81.118 67.645 ;
        RECT 76.012 64.225 84.462 64.301 ;
        RECT 81.072 59.165 81.118 67.645 ;
        RECT 72.608 67.629 81.072 67.691 ;
        RECT 76.058 64.179 84.508 64.255 ;
        RECT 81.026 59.211 81.072 67.691 ;
        RECT 72.562 67.675 81.026 67.737 ;
        RECT 76.104 64.133 84.554 64.209 ;
        RECT 80.98 59.257 81.026 67.737 ;
        RECT 72.516 67.721 80.98 67.783 ;
        RECT 76.15 64.087 84.6 64.163 ;
        RECT 80.934 59.303 80.98 67.783 ;
        RECT 72.47 67.767 80.934 67.829 ;
        RECT 76.196 64.041 84.646 64.117 ;
        RECT 80.888 59.349 80.934 67.829 ;
        RECT 72.424 67.813 80.888 67.875 ;
        RECT 76.242 63.995 84.692 64.071 ;
        RECT 80.842 59.395 80.888 67.875 ;
        RECT 72.378 67.859 80.842 67.921 ;
        RECT 76.288 63.949 84.738 64.025 ;
        RECT 80.796 59.441 80.842 67.921 ;
        RECT 72.332 67.905 80.796 67.967 ;
        RECT 76.334 63.903 84.784 63.979 ;
        RECT 80.75 59.487 80.796 67.967 ;
        RECT 72.286 67.951 80.75 68.013 ;
        RECT 76.38 63.857 84.83 63.933 ;
        RECT 80.704 59.533 80.75 68.013 ;
        RECT 72.24 67.997 80.704 68.059 ;
        RECT 76.426 63.811 84.876 63.887 ;
        RECT 80.658 59.579 80.704 68.059 ;
        RECT 72.194 68.043 80.658 68.105 ;
        RECT 76.472 63.765 84.922 63.841 ;
        RECT 80.612 59.625 80.658 68.105 ;
        RECT 72.148 68.089 80.612 68.151 ;
        RECT 76.518 63.719 84.968 63.795 ;
        RECT 80.566 59.671 80.612 68.151 ;
        RECT 72.102 68.135 80.566 68.197 ;
        RECT 76.564 63.673 85.014 63.749 ;
        RECT 80.52 59.717 80.566 68.197 ;
        RECT 72.056 68.181 80.52 68.243 ;
        RECT 76.61 63.627 85.06 63.703 ;
        RECT 80.474 59.763 80.52 68.243 ;
        RECT 72.01 68.227 80.474 68.289 ;
        RECT 76.656 63.581 85.106 63.657 ;
        RECT 80.428 59.809 80.474 68.289 ;
        RECT 71.964 68.273 80.428 68.335 ;
        RECT 76.702 63.535 85.152 63.611 ;
        RECT 80.382 59.855 80.428 68.335 ;
        RECT 71.918 68.319 80.382 68.381 ;
        RECT 76.748 63.489 85.198 63.565 ;
        RECT 80.336 59.901 80.382 68.381 ;
        RECT 71.872 68.365 80.336 68.427 ;
        RECT 76.794 63.443 110 63.5 ;
        RECT 80.29 59.947 80.336 68.427 ;
        RECT 71.826 68.411 80.29 68.473 ;
        RECT 76.84 63.397 110 63.5 ;
        RECT 80.244 59.993 80.29 68.473 ;
        RECT 71.78 68.457 80.244 68.519 ;
        RECT 76.886 63.351 110 63.5 ;
        RECT 80.198 60.039 80.244 68.519 ;
        RECT 71.734 68.503 80.198 68.565 ;
        RECT 76.932 63.305 110 63.5 ;
        RECT 80.152 60.085 80.198 68.565 ;
        RECT 71.688 68.549 80.152 68.611 ;
        RECT 76.978 63.259 110 63.5 ;
        RECT 80.106 60.131 80.152 68.611 ;
        RECT 71.642 68.595 80.106 68.657 ;
        RECT 77.024 63.213 110 63.5 ;
        RECT 80.06 60.177 80.106 68.657 ;
        RECT 71.596 68.641 80.06 68.703 ;
        RECT 77.07 63.167 110 63.5 ;
        RECT 80.014 60.223 80.06 68.703 ;
        RECT 71.55 68.687 80.014 68.749 ;
        RECT 77.116 63.121 110 63.5 ;
        RECT 79.968 60.269 80.014 68.749 ;
        RECT 71.504 68.733 79.968 68.795 ;
        RECT 77.162 63.075 110 63.5 ;
        RECT 79.922 60.315 79.968 68.795 ;
        RECT 71.458 68.779 79.922 68.841 ;
        RECT 77.208 63.029 110 63.5 ;
        RECT 79.876 60.361 79.922 68.841 ;
        RECT 71.412 68.825 79.876 68.887 ;
        RECT 77.254 62.983 110 63.5 ;
        RECT 79.83 60.407 79.876 68.887 ;
        RECT 71.366 68.871 79.83 68.933 ;
        RECT 77.3 62.937 110 63.5 ;
        RECT 79.784 60.453 79.83 68.933 ;
        RECT 71.32 68.917 79.784 68.979 ;
        RECT 77.346 62.891 110 63.5 ;
        RECT 79.738 60.499 79.784 68.979 ;
        RECT 71.274 68.963 79.738 69.025 ;
        RECT 77.392 62.845 110 63.5 ;
        RECT 79.692 60.545 79.738 69.025 ;
        RECT 71.228 69.009 79.692 69.071 ;
        RECT 77.438 62.799 110 63.5 ;
        RECT 79.646 60.591 79.692 69.071 ;
        RECT 71.182 69.055 79.646 69.117 ;
        RECT 77.484 62.753 110 63.5 ;
        RECT 79.6 60.637 79.646 69.117 ;
        RECT 71.136 69.101 79.6 69.163 ;
        RECT 77.53 62.707 110 63.5 ;
        RECT 79.554 60.683 79.6 69.163 ;
        RECT 71.09 69.147 79.554 69.209 ;
        RECT 77.576 62.661 110 63.5 ;
        RECT 79.508 60.729 79.554 69.209 ;
        RECT 71.044 69.193 79.508 69.255 ;
        RECT 77.622 62.615 110 63.5 ;
        RECT 79.462 60.775 79.508 69.255 ;
        RECT 70.998 69.239 79.462 69.301 ;
        RECT 77.668 62.569 110 63.5 ;
        RECT 79.416 60.821 79.462 69.301 ;
        RECT 70.952 69.285 79.416 69.347 ;
        RECT 77.714 62.523 110 63.5 ;
        RECT 79.37 60.867 79.416 69.347 ;
        RECT 70.906 69.331 79.37 69.393 ;
        RECT 77.76 62.477 110 63.5 ;
        RECT 79.324 60.913 79.37 69.393 ;
        RECT 70.86 69.377 79.324 69.439 ;
        RECT 77.806 62.431 110 63.5 ;
        RECT 79.278 60.959 79.324 69.439 ;
        RECT 69.515 30.5 110 42.5 ;
        RECT 57.496 42.496 74.483 42.524 ;
        RECT 52.574 47.418 69.515 47.477 ;
        RECT 52.62 47.372 69.561 47.447 ;
        RECT 69.502 30.506 69.515 47.477 ;
        RECT 52.666 47.326 69.607 47.401 ;
        RECT 69.456 30.536 69.502 47.506 ;
        RECT 52.528 47.464 69.456 47.552 ;
        RECT 52.712 47.28 69.653 47.355 ;
        RECT 69.41 30.582 69.456 47.552 ;
        RECT 52.482 47.51 69.41 47.598 ;
        RECT 52.758 47.234 69.699 47.309 ;
        RECT 69.364 30.628 69.41 47.598 ;
        RECT 52.436 47.556 69.364 47.644 ;
        RECT 52.804 47.188 69.745 47.263 ;
        RECT 69.318 30.674 69.364 47.644 ;
        RECT 52.39 47.602 69.318 47.69 ;
        RECT 52.85 47.142 69.791 47.217 ;
        RECT 69.272 30.72 69.318 47.69 ;
        RECT 52.344 47.648 69.272 47.736 ;
        RECT 52.896 47.096 69.837 47.171 ;
        RECT 69.226 30.766 69.272 47.736 ;
        RECT 52.298 47.694 69.226 47.782 ;
        RECT 52.942 47.05 69.883 47.125 ;
        RECT 69.18 30.812 69.226 47.782 ;
        RECT 52.252 47.74 69.18 47.828 ;
        RECT 52.988 47.004 69.929 47.079 ;
        RECT 69.134 30.858 69.18 47.828 ;
        RECT 52.206 47.786 69.134 47.874 ;
        RECT 53.034 46.958 69.975 47.033 ;
        RECT 69.088 30.904 69.134 47.874 ;
        RECT 52.16 47.832 69.088 47.92 ;
        RECT 53.08 46.912 70.021 46.987 ;
        RECT 69.042 30.95 69.088 47.92 ;
        RECT 52.114 47.878 69.042 47.966 ;
        RECT 53.126 46.866 70.067 46.941 ;
        RECT 68.996 30.996 69.042 47.966 ;
        RECT 52.068 47.924 68.996 48.012 ;
        RECT 53.172 46.82 70.113 46.895 ;
        RECT 68.95 31.042 68.996 48.012 ;
        RECT 52.022 47.97 68.95 48.058 ;
        RECT 53.218 46.774 70.159 46.849 ;
        RECT 68.904 31.088 68.95 48.058 ;
        RECT 51.976 48.016 68.904 48.104 ;
        RECT 53.264 46.728 70.205 46.803 ;
        RECT 68.858 31.134 68.904 48.104 ;
        RECT 51.93 48.062 68.858 48.15 ;
        RECT 53.31 46.682 70.251 46.757 ;
        RECT 68.812 31.18 68.858 48.15 ;
        RECT 51.884 48.108 68.812 48.196 ;
        RECT 53.356 46.636 70.297 46.711 ;
        RECT 68.766 31.226 68.812 48.196 ;
        RECT 51.838 48.154 68.766 48.242 ;
        RECT 53.402 46.59 70.343 46.665 ;
        RECT 68.72 31.272 68.766 48.242 ;
        RECT 51.792 48.2 68.72 48.288 ;
        RECT 53.448 46.544 70.389 46.619 ;
        RECT 68.674 31.318 68.72 48.288 ;
        RECT 51.746 48.246 68.674 48.334 ;
        RECT 53.494 46.498 70.435 46.573 ;
        RECT 68.628 31.364 68.674 48.334 ;
        RECT 51.7 48.292 68.628 48.38 ;
        RECT 53.54 46.452 70.481 46.527 ;
        RECT 68.582 31.41 68.628 48.38 ;
        RECT 51.654 48.338 68.582 48.426 ;
        RECT 53.586 46.406 70.527 46.481 ;
        RECT 68.536 31.456 68.582 48.426 ;
        RECT 51.608 48.384 68.536 48.472 ;
        RECT 53.632 46.36 70.573 46.435 ;
        RECT 68.49 31.502 68.536 48.472 ;
        RECT 51.562 48.43 68.49 48.518 ;
        RECT 53.678 46.314 70.619 46.389 ;
        RECT 68.444 31.548 68.49 48.518 ;
        RECT 51.516 48.476 68.444 48.564 ;
        RECT 53.724 46.268 70.665 46.343 ;
        RECT 68.398 31.594 68.444 48.564 ;
        RECT 51.47 48.522 68.398 48.61 ;
        RECT 53.77 46.222 70.711 46.297 ;
        RECT 68.352 31.64 68.398 48.61 ;
        RECT 51.424 48.568 68.352 48.656 ;
        RECT 53.816 46.176 70.757 46.251 ;
        RECT 68.306 31.686 68.352 48.656 ;
        RECT 51.378 48.614 68.306 48.702 ;
        RECT 53.862 46.13 70.803 46.205 ;
        RECT 68.26 31.732 68.306 48.702 ;
        RECT 51.332 48.66 68.26 48.748 ;
        RECT 53.908 46.084 70.849 46.159 ;
        RECT 68.214 31.778 68.26 48.748 ;
        RECT 51.286 48.706 68.214 48.794 ;
        RECT 53.954 46.038 70.895 46.113 ;
        RECT 68.168 31.824 68.214 48.794 ;
        RECT 51.24 48.752 68.168 48.84 ;
        RECT 54 45.992 70.941 46.067 ;
        RECT 68.122 31.87 68.168 48.84 ;
        RECT 51.194 48.798 68.122 48.886 ;
        RECT 54.046 45.946 70.987 46.021 ;
        RECT 68.076 31.916 68.122 48.886 ;
        RECT 51.148 48.844 68.076 48.932 ;
        RECT 54.092 45.9 71.033 45.975 ;
        RECT 68.03 31.962 68.076 48.932 ;
        RECT 51.102 48.89 68.03 48.978 ;
        RECT 54.138 45.854 71.079 45.929 ;
        RECT 67.984 32.008 68.03 48.978 ;
        RECT 51.056 48.936 67.984 49.024 ;
        RECT 54.184 45.808 71.125 45.883 ;
        RECT 67.938 32.054 67.984 49.024 ;
        RECT 51.01 48.982 67.938 49.07 ;
        RECT 54.23 45.762 71.171 45.837 ;
        RECT 67.892 32.1 67.938 49.07 ;
        RECT 50.964 49.028 67.892 49.116 ;
        RECT 54.276 45.716 71.217 45.791 ;
        RECT 67.846 32.146 67.892 49.116 ;
        RECT 50.918 49.074 67.846 49.162 ;
        RECT 54.322 45.67 71.263 45.745 ;
        RECT 67.8 32.192 67.846 49.162 ;
        RECT 50.872 49.12 67.8 49.208 ;
        RECT 54.368 45.624 71.309 45.699 ;
        RECT 67.754 32.238 67.8 49.208 ;
        RECT 50.826 49.166 67.754 49.254 ;
        RECT 54.414 45.578 71.355 45.653 ;
        RECT 67.708 32.284 67.754 49.254 ;
        RECT 50.78 49.212 67.708 49.3 ;
        RECT 54.46 45.532 71.401 45.607 ;
        RECT 67.662 32.33 67.708 49.3 ;
        RECT 50.734 49.258 67.662 49.346 ;
        RECT 54.506 45.486 71.447 45.561 ;
        RECT 67.616 32.376 67.662 49.346 ;
        RECT 50.688 49.304 67.616 49.392 ;
        RECT 54.552 45.44 71.493 45.515 ;
        RECT 67.57 32.422 67.616 49.392 ;
        RECT 50.642 49.35 67.57 49.438 ;
        RECT 54.598 45.394 71.539 45.469 ;
        RECT 67.524 32.468 67.57 49.438 ;
        RECT 50.596 49.396 67.524 49.484 ;
        RECT 54.644 45.348 71.585 45.423 ;
        RECT 67.478 32.514 67.524 49.484 ;
        RECT 50.55 49.442 67.478 49.53 ;
        RECT 54.69 45.302 71.631 45.377 ;
        RECT 67.432 32.56 67.478 49.53 ;
        RECT 50.504 49.488 67.432 49.576 ;
        RECT 54.736 45.256 71.677 45.331 ;
        RECT 67.386 32.606 67.432 49.576 ;
        RECT 50.458 49.534 67.386 49.622 ;
        RECT 54.782 45.21 71.723 45.285 ;
        RECT 67.34 32.652 67.386 49.622 ;
        RECT 50.412 49.58 67.34 49.668 ;
        RECT 54.828 45.164 71.769 45.239 ;
        RECT 67.294 32.698 67.34 49.668 ;
        RECT 50.366 49.626 67.294 49.714 ;
        RECT 54.874 45.118 71.815 45.193 ;
        RECT 67.248 32.744 67.294 49.714 ;
        RECT 50.32 49.672 67.248 49.76 ;
        RECT 54.92 45.072 71.861 45.147 ;
        RECT 67.202 32.79 67.248 49.76 ;
        RECT 50.274 49.718 67.202 49.806 ;
        RECT 54.966 45.026 71.907 45.101 ;
        RECT 67.156 32.836 67.202 49.806 ;
        RECT 50.228 49.764 67.156 49.852 ;
        RECT 55.012 44.98 71.953 45.055 ;
        RECT 67.11 32.882 67.156 49.852 ;
        RECT 50.182 49.81 67.11 49.898 ;
        RECT 55.058 44.934 71.999 45.009 ;
        RECT 67.064 32.928 67.11 49.898 ;
        RECT 50.136 49.856 67.064 49.944 ;
        RECT 55.104 44.888 72.045 44.963 ;
        RECT 67.018 32.974 67.064 49.944 ;
        RECT 50.09 49.902 67.018 49.99 ;
        RECT 55.15 44.842 72.091 44.917 ;
        RECT 66.972 33.02 67.018 49.99 ;
        RECT 50.044 49.948 66.972 50.036 ;
        RECT 55.196 44.796 72.137 44.871 ;
        RECT 66.926 33.066 66.972 50.036 ;
        RECT 49.998 49.994 66.926 50.082 ;
        RECT 55.242 44.75 72.183 44.825 ;
        RECT 66.88 33.112 66.926 50.082 ;
        RECT 49.952 50.04 66.88 50.128 ;
        RECT 55.288 44.704 72.229 44.779 ;
        RECT 66.834 33.158 66.88 50.128 ;
        RECT 49.906 50.086 66.834 50.174 ;
        RECT 55.334 44.658 72.275 44.733 ;
        RECT 66.788 33.204 66.834 50.174 ;
        RECT 49.86 50.132 66.788 50.22 ;
        RECT 55.38 44.612 72.321 44.687 ;
        RECT 66.742 33.25 66.788 50.22 ;
        RECT 49.814 50.178 66.742 50.266 ;
        RECT 55.426 44.566 72.367 44.641 ;
        RECT 66.696 33.296 66.742 50.266 ;
        RECT 49.768 50.224 66.696 50.312 ;
        RECT 55.472 44.52 72.413 44.595 ;
        RECT 66.65 33.342 66.696 50.312 ;
        RECT 49.722 50.27 66.65 50.358 ;
        RECT 55.518 44.474 72.459 44.549 ;
        RECT 66.604 33.388 66.65 50.358 ;
        RECT 49.676 50.316 66.604 50.404 ;
        RECT 55.564 44.428 72.505 44.503 ;
        RECT 66.558 33.434 66.604 50.404 ;
        RECT 49.63 50.362 66.558 50.45 ;
        RECT 55.61 44.382 72.551 44.457 ;
        RECT 66.512 33.48 66.558 50.45 ;
        RECT 49.584 50.408 66.512 50.496 ;
        RECT 55.656 44.336 72.597 44.411 ;
        RECT 66.466 33.526 66.512 50.496 ;
        RECT 49.538 50.454 66.466 50.542 ;
        RECT 55.702 44.29 72.643 44.365 ;
        RECT 66.42 33.572 66.466 50.542 ;
        RECT 49.492 50.5 66.42 50.588 ;
        RECT 55.748 44.244 72.689 44.319 ;
        RECT 66.374 33.618 66.42 50.588 ;
        RECT 49.446 50.546 66.374 50.634 ;
        RECT 55.794 44.198 72.735 44.273 ;
        RECT 66.328 33.664 66.374 50.634 ;
        RECT 49.4 50.592 66.328 50.68 ;
        RECT 55.84 44.152 72.781 44.227 ;
        RECT 66.282 33.71 66.328 50.68 ;
        RECT 49.354 50.638 66.282 50.726 ;
        RECT 55.886 44.106 72.827 44.181 ;
        RECT 66.236 33.756 66.282 50.726 ;
        RECT 49.308 50.684 66.236 50.772 ;
        RECT 55.932 44.06 72.873 44.135 ;
        RECT 66.19 33.802 66.236 50.772 ;
        RECT 49.262 50.73 66.19 50.818 ;
        RECT 55.978 44.014 72.919 44.089 ;
        RECT 66.144 33.848 66.19 50.818 ;
        RECT 49.216 50.776 66.144 50.864 ;
        RECT 56.024 43.968 72.965 44.043 ;
        RECT 66.098 33.894 66.144 50.864 ;
        RECT 49.17 50.822 66.098 50.91 ;
        RECT 56.07 43.922 73.011 43.997 ;
        RECT 66.052 33.94 66.098 50.91 ;
        RECT 49.124 50.868 66.052 50.956 ;
        RECT 56.116 43.876 73.057 43.951 ;
        RECT 66.006 33.986 66.052 50.956 ;
        RECT 49.078 50.914 66.006 51.002 ;
        RECT 56.162 43.83 73.103 43.905 ;
        RECT 65.96 34.032 66.006 51.002 ;
        RECT 49.032 50.96 65.96 51.048 ;
        RECT 56.208 43.784 73.149 43.859 ;
        RECT 65.914 34.078 65.96 51.048 ;
        RECT 48.986 51.006 65.914 51.094 ;
        RECT 56.254 43.738 73.195 43.813 ;
        RECT 65.868 34.124 65.914 51.094 ;
        RECT 48.94 51.052 65.868 51.14 ;
        RECT 56.3 43.692 73.241 43.767 ;
        RECT 65.822 34.17 65.868 51.14 ;
        RECT 48.894 51.098 65.822 51.186 ;
        RECT 56.346 43.646 73.287 43.721 ;
        RECT 65.776 34.216 65.822 51.186 ;
        RECT 48.848 51.144 65.776 51.232 ;
        RECT 56.392 43.6 73.333 43.675 ;
        RECT 65.73 34.262 65.776 51.232 ;
        RECT 48.802 51.19 65.73 51.278 ;
        RECT 56.438 43.554 73.379 43.629 ;
        RECT 65.684 34.308 65.73 51.278 ;
        RECT 48.756 51.236 65.684 51.324 ;
        RECT 56.484 43.508 73.425 43.583 ;
        RECT 65.638 34.354 65.684 51.324 ;
        RECT 48.71 51.282 65.638 51.37 ;
        RECT 56.53 43.462 73.471 43.537 ;
        RECT 65.592 34.4 65.638 51.37 ;
        RECT 48.664 51.328 65.592 51.416 ;
        RECT 56.576 43.416 73.517 43.491 ;
        RECT 65.546 34.446 65.592 51.416 ;
        RECT 48.618 51.374 65.546 51.462 ;
        RECT 56.622 43.37 73.563 43.445 ;
        RECT 65.5 34.492 65.546 51.462 ;
        RECT 48.572 51.42 65.5 51.508 ;
        RECT 56.668 43.324 73.609 43.399 ;
        RECT 65.454 34.538 65.5 51.508 ;
        RECT 48.526 51.466 65.454 51.554 ;
        RECT 56.714 43.278 73.655 43.353 ;
        RECT 65.408 34.584 65.454 51.554 ;
        RECT 48.48 51.512 65.408 51.6 ;
        RECT 56.76 43.232 73.701 43.307 ;
        RECT 65.362 34.63 65.408 51.6 ;
        RECT 48.434 51.558 65.362 51.646 ;
        RECT 56.806 43.186 73.747 43.261 ;
        RECT 65.316 34.676 65.362 51.646 ;
        RECT 48.388 51.604 65.316 51.692 ;
        RECT 56.852 43.14 73.793 43.215 ;
        RECT 65.27 34.722 65.316 51.692 ;
        RECT 48.342 51.65 65.27 51.738 ;
        RECT 56.898 43.094 73.839 43.169 ;
        RECT 65.224 34.768 65.27 51.738 ;
        RECT 48.296 51.696 65.224 51.784 ;
        RECT 56.944 43.048 73.885 43.123 ;
        RECT 65.178 34.814 65.224 51.784 ;
        RECT 48.25 51.742 65.178 51.83 ;
        RECT 56.99 43.002 73.931 43.077 ;
        RECT 65.132 34.86 65.178 51.83 ;
        RECT 48.204 51.788 65.132 51.876 ;
        RECT 57.036 42.956 73.977 43.031 ;
        RECT 65.086 34.906 65.132 51.876 ;
        RECT 48.158 51.834 65.086 51.922 ;
        RECT 57.082 42.91 74.023 42.985 ;
        RECT 65.04 34.952 65.086 51.922 ;
        RECT 48.112 51.88 65.04 51.968 ;
        RECT 57.128 42.864 74.069 42.939 ;
        RECT 64.994 34.998 65.04 51.968 ;
        RECT 48.066 51.926 64.994 52.014 ;
        RECT 57.174 42.818 74.115 42.893 ;
        RECT 64.948 35.044 64.994 52.014 ;
        RECT 48.02 51.972 64.948 52.06 ;
        RECT 57.22 42.772 74.161 42.847 ;
        RECT 64.902 35.09 64.948 52.06 ;
        RECT 47.974 52.018 64.902 52.106 ;
        RECT 57.266 42.726 74.207 42.801 ;
        RECT 64.856 35.136 64.902 52.106 ;
        RECT 47.928 52.064 64.856 52.152 ;
        RECT 57.312 42.68 74.253 42.755 ;
        RECT 64.81 35.182 64.856 52.152 ;
        RECT 47.882 52.11 64.81 52.198 ;
        RECT 57.358 42.634 74.299 42.709 ;
        RECT 64.764 35.228 64.81 52.198 ;
        RECT 47.836 52.156 64.764 52.244 ;
        RECT 57.404 42.588 74.345 42.663 ;
        RECT 64.718 35.274 64.764 52.244 ;
        RECT 47.79 52.202 64.718 52.29 ;
        RECT 57.45 42.542 74.391 42.617 ;
        RECT 64.672 35.32 64.718 52.29 ;
        RECT 47.744 52.248 64.672 52.336 ;
        RECT 57.496 42.496 74.437 42.571 ;
        RECT 64.626 35.366 64.672 52.336 ;
        RECT 47.698 52.294 64.626 52.382 ;
        RECT 57.542 42.45 110 42.5 ;
        RECT 64.58 35.412 64.626 52.382 ;
        RECT 47.652 52.34 64.58 52.428 ;
        RECT 57.588 42.404 110 42.5 ;
        RECT 64.534 35.458 64.58 52.428 ;
        RECT 47.606 52.386 64.534 52.474 ;
        RECT 57.634 42.358 110 42.5 ;
        RECT 64.488 35.504 64.534 52.474 ;
        RECT 47.56 52.432 64.488 52.52 ;
        RECT 57.68 42.312 110 42.5 ;
        RECT 64.442 35.55 64.488 52.52 ;
        RECT 47.514 52.478 64.442 52.566 ;
        RECT 57.726 42.266 110 42.5 ;
        RECT 64.396 35.596 64.442 52.566 ;
        RECT 47.468 52.524 64.396 52.612 ;
        RECT 57.772 42.22 110 42.5 ;
        RECT 64.35 35.642 64.396 52.612 ;
        RECT 47.422 52.57 64.35 52.658 ;
        RECT 57.818 42.174 110 42.5 ;
        RECT 64.304 35.688 64.35 52.658 ;
        RECT 47.376 52.616 64.304 52.704 ;
        RECT 57.864 42.128 110 42.5 ;
        RECT 64.258 35.734 64.304 52.704 ;
        RECT 47.33 52.662 64.258 52.75 ;
        RECT 57.91 42.082 110 42.5 ;
        RECT 64.212 35.78 64.258 52.75 ;
        RECT 47.284 52.708 64.212 52.796 ;
        RECT 57.956 42.036 110 42.5 ;
        RECT 64.166 35.826 64.212 52.796 ;
        RECT 47.238 52.754 64.166 52.842 ;
        RECT 58.002 41.99 110 42.5 ;
        RECT 64.12 35.872 64.166 52.842 ;
        RECT 47.192 52.8 64.12 52.888 ;
        RECT 58.048 41.944 110 42.5 ;
        RECT 64.074 35.918 64.12 52.888 ;
        RECT 47.146 52.846 64.074 52.934 ;
        RECT 58.094 41.898 110 42.5 ;
        RECT 64.028 35.964 64.074 52.934 ;
        RECT 47.1 52.892 64.028 52.98 ;
        RECT 58.14 41.852 110 42.5 ;
        RECT 63.982 36.01 64.028 52.98 ;
        RECT 47.054 52.938 63.982 53.026 ;
        RECT 58.186 41.806 110 42.5 ;
        RECT 63.936 36.056 63.982 53.026 ;
        RECT 47.008 52.984 63.936 53.072 ;
        RECT 58.232 41.76 110 42.5 ;
        RECT 63.89 36.102 63.936 53.072 ;
        RECT 46.962 53.03 63.89 53.118 ;
        RECT 58.278 41.714 110 42.5 ;
        RECT 63.844 36.148 63.89 53.118 ;
        RECT 46.916 53.076 63.844 53.164 ;
        RECT 58.324 41.668 110 42.5 ;
        RECT 63.798 36.194 63.844 53.164 ;
        RECT 46.87 53.122 63.798 53.21 ;
        RECT 58.37 41.622 110 42.5 ;
        RECT 63.752 36.24 63.798 53.21 ;
        RECT 46.824 53.168 63.752 53.256 ;
        RECT 58.416 41.576 110 42.5 ;
        RECT 63.706 36.286 63.752 53.256 ;
        RECT 46.778 53.214 63.706 53.302 ;
        RECT 58.462 41.53 110 42.5 ;
        RECT 63.66 36.332 63.706 53.302 ;
        RECT 46.732 53.26 63.66 53.348 ;
        RECT 58.508 41.484 110 42.5 ;
        RECT 63.614 36.378 63.66 53.348 ;
        RECT 46.686 53.306 63.614 53.394 ;
        RECT 58.554 41.438 110 42.5 ;
        RECT 63.568 36.424 63.614 53.394 ;
        RECT 46.64 53.352 63.568 53.44 ;
        RECT 58.6 41.392 110 42.5 ;
        RECT 63.522 36.47 63.568 53.44 ;
        RECT 46.594 53.398 63.522 53.486 ;
        RECT 58.646 41.346 110 42.5 ;
        RECT 63.476 36.516 63.522 53.486 ;
        RECT 46.548 53.444 63.476 53.532 ;
        RECT 58.692 41.3 110 42.5 ;
        RECT 63.43 36.562 63.476 53.532 ;
        RECT 46.502 53.49 63.43 53.578 ;
        RECT 58.738 41.254 110 42.5 ;
        RECT 63.384 36.608 63.43 53.578 ;
        RECT 46.456 53.536 63.384 53.624 ;
        RECT 58.784 41.208 110 42.5 ;
        RECT 63.338 36.654 63.384 53.624 ;
        RECT 46.41 53.582 63.338 53.67 ;
        RECT 58.83 41.162 110 42.5 ;
        RECT 63.292 36.7 63.338 53.67 ;
        RECT 46.364 53.628 63.292 53.716 ;
        RECT 58.876 41.116 110 42.5 ;
        RECT 63.246 36.746 63.292 53.716 ;
        RECT 46.318 53.674 63.246 53.762 ;
        RECT 58.922 41.07 110 42.5 ;
        RECT 63.2 36.792 63.246 53.762 ;
        RECT 46.272 53.72 63.2 53.808 ;
        RECT 58.968 41.024 110 42.5 ;
        RECT 63.154 36.838 63.2 53.808 ;
        RECT 46.226 53.766 63.154 53.854 ;
        RECT 59.014 40.978 110 42.5 ;
        RECT 63.108 36.884 63.154 53.854 ;
        RECT 46.18 53.812 63.108 53.9 ;
        RECT 59.06 40.932 110 42.5 ;
        RECT 63.062 36.93 63.108 53.9 ;
        RECT 46.134 53.858 63.062 53.946 ;
        RECT 59.106 40.886 110 42.5 ;
        RECT 63.016 36.976 63.062 53.946 ;
        RECT 46.088 53.904 63.016 53.992 ;
        RECT 59.152 40.84 110 42.5 ;
        RECT 62.97 37.022 63.016 53.992 ;
        RECT 46.042 53.95 62.97 54.038 ;
        RECT 59.198 40.794 110 42.5 ;
        RECT 62.924 37.068 62.97 54.038 ;
        RECT 45.996 53.996 62.924 54.084 ;
        RECT 59.244 40.748 110 42.5 ;
        RECT 62.878 37.114 62.924 54.084 ;
        RECT 45.95 54.042 62.878 54.13 ;
        RECT 59.29 40.702 110 42.5 ;
        RECT 62.832 37.16 62.878 54.13 ;
        RECT 45.904 54.088 62.832 54.176 ;
        RECT 59.336 40.656 110 42.5 ;
        RECT 62.786 37.206 62.832 54.176 ;
        RECT 45.858 54.134 62.786 54.222 ;
        RECT 59.382 40.61 110 42.5 ;
        RECT 62.74 37.252 62.786 54.222 ;
        RECT 45.812 54.18 62.74 54.268 ;
        RECT 59.428 40.564 110 42.5 ;
        RECT 62.694 37.298 62.74 54.268 ;
        RECT 45.766 54.226 62.694 54.314 ;
        RECT 59.474 40.518 110 42.5 ;
        RECT 62.648 37.344 62.694 54.314 ;
        RECT 45.72 54.272 62.648 54.36 ;
        RECT 59.52 40.472 110 42.5 ;
        RECT 62.602 37.39 62.648 54.36 ;
        RECT 45.674 54.318 62.602 54.406 ;
        RECT 59.566 40.426 110 42.5 ;
        RECT 62.556 37.436 62.602 54.406 ;
        RECT 45.628 54.364 62.556 54.452 ;
        RECT 59.612 40.38 110 42.5 ;
        RECT 62.51 37.482 62.556 54.452 ;
        RECT 45.582 54.41 62.51 54.498 ;
        RECT 59.658 40.334 110 42.5 ;
        RECT 62.464 37.528 62.51 54.498 ;
        RECT 45.536 54.456 62.464 54.544 ;
        RECT 59.704 40.288 110 42.5 ;
        RECT 62.418 37.574 62.464 54.544 ;
        RECT 45.49 54.502 62.418 54.59 ;
        RECT 59.75 40.242 110 42.5 ;
        RECT 62.372 37.62 62.418 54.59 ;
        RECT 45.444 54.548 62.372 54.636 ;
        RECT 59.796 40.196 110 42.5 ;
        RECT 62.326 37.666 62.372 54.636 ;
        RECT 45.398 54.594 62.326 54.682 ;
        RECT 59.842 40.15 110 42.5 ;
        RECT 62.28 37.712 62.326 54.682 ;
        RECT 45.352 54.64 62.28 54.728 ;
        RECT 59.888 40.104 110 42.5 ;
        RECT 62.234 37.758 62.28 54.728 ;
        RECT 45.306 54.686 62.234 54.774 ;
        RECT 59.934 40.058 110 42.5 ;
        RECT 62.188 37.804 62.234 54.774 ;
        RECT 45.26 54.732 62.188 54.82 ;
        RECT 59.98 40.012 110 42.5 ;
        RECT 62.142 37.85 62.188 54.82 ;
        RECT 45.214 54.778 62.142 54.866 ;
        RECT 60.026 39.966 110 42.5 ;
        RECT 62.096 37.896 62.142 54.866 ;
        RECT 45.168 54.824 62.096 54.912 ;
        RECT 60.072 39.92 110 42.5 ;
        RECT 62.05 37.942 62.096 54.912 ;
        RECT 45.122 54.87 62.05 54.958 ;
        RECT 60.118 39.874 110 42.5 ;
        RECT 62.004 37.988 62.05 54.958 ;
        RECT 45.076 54.916 62.004 55.004 ;
        RECT 60.164 39.828 110 42.5 ;
        RECT 61.958 38.034 62.004 55.004 ;
        RECT 45.03 54.962 61.958 55.05 ;
        RECT 60.21 39.782 110 42.5 ;
        RECT 61.912 38.08 61.958 55.05 ;
        RECT 44.984 55.008 61.912 55.096 ;
        RECT 60.256 39.736 110 42.5 ;
        RECT 61.866 38.126 61.912 55.096 ;
        RECT 44.938 55.054 61.866 55.142 ;
        RECT 60.302 39.69 110 42.5 ;
        RECT 61.82 38.172 61.866 55.142 ;
        RECT 44.892 55.1 61.82 55.188 ;
        RECT 60.348 39.644 110 42.5 ;
        RECT 61.774 38.218 61.82 55.188 ;
        RECT 44.846 55.146 61.774 55.234 ;
        RECT 60.394 39.598 110 42.5 ;
        RECT 61.728 38.264 61.774 55.234 ;
        RECT 44.8 55.192 61.728 55.28 ;
        RECT 60.44 39.552 110 42.5 ;
        RECT 61.682 38.31 61.728 55.28 ;
        RECT 44.754 55.238 61.682 55.326 ;
        RECT 60.486 39.506 110 42.5 ;
        RECT 61.636 38.356 61.682 55.326 ;
        RECT 44.708 55.284 61.636 55.372 ;
        RECT 60.532 39.46 110 42.5 ;
        RECT 61.59 38.402 61.636 55.372 ;
        RECT 44.662 55.33 61.59 55.418 ;
        RECT 60.578 39.414 110 42.5 ;
        RECT 61.544 38.448 61.59 55.418 ;
        RECT 44.616 55.376 61.544 55.464 ;
        RECT 60.624 39.368 110 42.5 ;
        RECT 61.498 38.494 61.544 55.464 ;
        RECT 44.57 55.422 61.498 55.51 ;
        RECT 60.67 39.322 110 42.5 ;
        RECT 61.452 38.54 61.498 55.51 ;
        RECT 44.524 55.468 61.452 55.556 ;
        RECT 60.716 39.276 110 42.5 ;
        RECT 61.406 38.586 61.452 55.556 ;
        RECT 44.478 55.514 61.406 55.602 ;
        RECT 60.762 39.23 110 42.5 ;
        RECT 61.36 38.632 61.406 55.602 ;
        RECT 44.432 55.56 61.36 55.648 ;
        RECT 60.808 39.184 110 42.5 ;
        RECT 61.314 38.678 61.36 55.648 ;
        RECT 44.386 55.606 61.314 55.694 ;
        RECT 60.854 39.138 110 42.5 ;
        RECT 61.268 38.724 61.314 55.694 ;
        RECT 44.34 55.652 61.268 55.74 ;
        RECT 60.9 39.092 110 42.5 ;
        RECT 61.222 38.77 61.268 55.74 ;
        RECT 44.294 55.698 61.222 55.786 ;
        RECT 60.946 39.046 110 42.5 ;
        RECT 61.176 38.816 61.222 55.786 ;
        RECT 44.248 55.744 61.176 55.832 ;
        RECT 60.992 39 110 42.5 ;
        RECT 61.13 38.862 61.176 55.832 ;
        RECT 44.202 55.79 61.13 55.878 ;
        RECT 61.038 38.954 110 42.5 ;
        RECT 61.084 38.908 61.13 55.878 ;
        RECT 44.156 55.836 61.084 55.924 ;
        RECT 44.11 55.882 61.038 55.97 ;
        RECT 44.064 55.928 60.992 56.016 ;
        RECT 44.018 55.974 60.946 56.062 ;
        RECT 43.972 56.02 60.9 56.108 ;
        RECT 43.926 56.066 60.854 56.154 ;
        RECT 43.88 56.112 60.808 56.2 ;
        RECT 43.834 56.158 60.762 56.246 ;
        RECT 43.788 56.204 60.716 56.292 ;
        RECT 43.742 56.25 60.67 56.338 ;
        RECT 43.696 56.296 60.624 56.384 ;
        RECT 43.65 56.342 60.578 56.43 ;
        RECT 43.604 56.388 60.532 56.476 ;
        RECT 43.558 56.434 60.486 56.522 ;
        RECT 43.512 56.48 60.44 56.568 ;
        RECT 43.466 56.526 60.394 56.614 ;
        RECT 43.42 56.572 60.348 56.66 ;
        RECT 43.374 56.618 60.302 56.706 ;
        RECT 43.328 56.664 60.256 56.752 ;
        RECT 43.282 56.71 60.21 56.798 ;
        RECT 43.236 56.756 60.164 56.844 ;
        RECT 43.19 56.802 60.118 56.89 ;
        RECT 43.144 56.848 60.072 56.936 ;
        RECT 43.098 56.894 60.026 56.982 ;
        RECT 43.052 56.94 59.98 57.028 ;
        RECT 43.006 56.986 59.934 57.074 ;
        RECT 42.96 57.032 59.888 57.12 ;
        RECT 42.914 57.078 59.842 57.166 ;
        RECT 42.868 57.124 59.796 57.212 ;
        RECT 42.822 57.17 59.75 57.258 ;
        RECT 42.776 57.216 59.704 57.304 ;
        RECT 42.73 57.262 59.658 57.35 ;
        RECT 42.684 57.308 59.612 57.396 ;
        RECT 42.638 57.354 59.566 57.442 ;
        RECT 42.592 57.4 59.52 57.488 ;
        RECT 42.5 57.492 59.474 57.534 ;
        RECT 42.546 57.446 59.474 57.534 ;
        RECT 42.46 57.535 59.428 57.58 ;
        RECT 42.414 57.578 59.382 57.626 ;
        RECT 42.368 57.624 59.336 57.672 ;
        RECT 42.322 57.67 59.29 57.718 ;
        RECT 42.276 57.716 59.244 57.764 ;
        RECT 42.23 57.762 59.198 57.81 ;
        RECT 42.184 57.808 59.152 57.856 ;
        RECT 42.138 57.854 59.106 57.902 ;
        RECT 42.092 57.9 59.06 57.948 ;
        RECT 42.046 57.946 59.014 57.994 ;
        RECT 42 57.992 58.968 58.04 ;
        RECT 41.954 58.038 58.922 58.086 ;
        RECT 41.908 58.084 58.876 58.132 ;
        RECT 41.862 58.13 58.83 58.178 ;
        RECT 41.816 58.176 58.784 58.224 ;
        RECT 41.77 58.222 58.738 58.27 ;
        RECT 41.724 58.268 58.692 58.316 ;
        RECT 41.678 58.314 58.646 58.362 ;
        RECT 41.632 58.36 58.6 58.408 ;
        RECT 41.586 58.406 58.554 58.454 ;
        RECT 41.54 58.452 58.508 58.5 ;
        RECT 41.494 58.498 58.462 58.546 ;
        RECT 41.448 58.544 58.416 58.592 ;
        RECT 41.402 58.59 58.37 58.638 ;
        RECT 41.356 58.636 58.324 58.684 ;
        RECT 41.31 58.682 58.278 58.73 ;
        RECT 41.264 58.728 58.232 58.776 ;
        RECT 41.218 58.774 58.186 58.822 ;
        RECT 41.172 58.82 58.14 58.868 ;
        RECT 41.126 58.866 58.094 58.914 ;
        RECT 41.08 58.912 58.048 58.96 ;
        RECT 41.034 58.958 58.002 59.006 ;
        RECT 40.988 59.004 57.956 59.052 ;
        RECT 40.942 59.05 57.91 59.098 ;
        RECT 40.896 59.096 57.864 59.144 ;
        RECT 40.85 59.142 57.818 59.19 ;
        RECT 40.804 59.188 57.772 59.236 ;
        RECT 40.758 59.234 57.726 59.282 ;
        RECT 40.712 59.28 57.68 59.328 ;
        RECT 40.666 59.326 57.634 59.374 ;
        RECT 40.62 59.372 57.588 59.42 ;
        RECT 40.574 59.418 57.542 59.466 ;
        RECT 40.528 59.464 57.496 59.512 ;
        RECT 40.482 59.51 57.45 59.558 ;
        RECT 40.436 59.556 57.404 59.604 ;
        RECT 40.39 59.602 57.358 59.65 ;
        RECT 40.344 59.648 57.312 59.696 ;
        RECT 40.298 59.694 57.266 59.742 ;
        RECT 40.252 59.74 57.22 59.788 ;
        RECT 40.206 59.786 57.174 59.834 ;
        RECT 40.16 59.832 57.128 59.88 ;
        RECT 40.114 59.878 57.082 59.926 ;
        RECT 40.068 59.924 57.036 59.972 ;
        RECT 40.022 59.97 56.99 60.018 ;
        RECT 39.976 60.016 56.944 60.064 ;
        RECT 39.93 60.062 56.898 60.11 ;
        RECT 39.884 60.108 56.852 60.156 ;
        RECT 39.838 60.154 56.806 60.202 ;
        RECT 39.792 60.2 56.76 60.248 ;
        RECT 39.746 60.246 56.714 60.294 ;
        RECT 39.7 60.292 56.668 60.34 ;
        RECT 39.654 60.338 56.622 60.386 ;
        RECT 39.608 60.384 56.576 60.432 ;
        RECT 39.562 60.43 56.53 60.478 ;
        RECT 39.516 60.476 56.484 60.524 ;
        RECT 39.47 60.522 56.438 60.57 ;
        RECT 39.424 60.568 56.392 60.616 ;
        RECT 39.378 60.614 56.346 60.662 ;
        RECT 39.332 60.66 56.3 60.708 ;
        RECT 39.286 60.706 56.254 60.754 ;
        RECT 39.24 60.752 56.208 60.8 ;
        RECT 39.194 60.798 56.162 60.846 ;
        RECT 39.148 60.844 56.116 60.892 ;
        RECT 39.102 60.89 56.07 60.938 ;
        RECT 39.056 60.936 56.024 60.984 ;
        RECT 39.01 60.982 55.978 61.03 ;
        RECT 38.964 61.028 55.932 61.076 ;
        RECT 38.918 61.074 55.886 61.122 ;
        RECT 38.872 61.12 55.84 61.168 ;
        RECT 38.826 61.166 55.794 61.214 ;
        RECT 38.78 61.212 55.748 61.26 ;
        RECT 38.734 61.258 55.702 61.306 ;
        RECT 38.688 61.304 55.656 61.352 ;
        RECT 38.642 61.35 55.61 61.398 ;
        RECT 38.596 61.396 55.564 61.444 ;
        RECT 38.55 61.442 55.518 61.49 ;
        RECT 38.504 61.488 55.472 61.536 ;
        RECT 38.458 61.534 55.426 61.582 ;
        RECT 38.412 61.58 55.38 61.628 ;
        RECT 38.366 61.626 55.334 61.674 ;
        RECT 38.32 61.672 55.288 61.72 ;
        RECT 38.274 61.718 55.242 61.766 ;
        RECT 38.228 61.764 55.196 61.812 ;
        RECT 38.182 61.81 55.15 61.858 ;
        RECT 38.136 61.856 55.104 61.904 ;
        RECT 38.09 61.902 55.058 61.95 ;
        RECT 38.044 61.948 55.012 61.996 ;
        RECT 37.998 61.994 54.966 62.042 ;
        RECT 37.952 62.04 54.92 62.088 ;
        RECT 37.906 62.086 54.874 62.134 ;
        RECT 37.86 62.132 54.828 62.18 ;
        RECT 37.814 62.178 54.782 62.226 ;
        RECT 37.768 62.224 54.736 62.272 ;
        RECT 37.722 62.27 54.69 62.318 ;
        RECT 37.676 62.316 54.644 62.364 ;
        RECT 37.63 62.362 54.598 62.41 ;
        RECT 37.584 62.408 54.552 62.456 ;
        RECT 37.538 62.454 54.506 62.502 ;
        RECT 37.492 62.5 54.46 62.548 ;
        RECT 37.446 62.546 54.414 62.594 ;
        RECT 37.4 62.592 54.368 62.64 ;
        RECT 37.354 62.638 54.322 62.686 ;
        RECT 37.308 62.684 54.276 62.732 ;
        RECT 37.262 62.73 54.23 62.778 ;
        RECT 37.216 62.776 54.184 62.824 ;
        RECT 37.17 62.822 54.138 62.87 ;
        RECT 37.124 62.868 54.092 62.916 ;
        RECT 37.078 62.914 54.046 62.962 ;
        RECT 37.032 62.96 54 63.008 ;
        RECT 36.986 63.006 53.954 63.054 ;
        RECT 36.94 63.052 53.908 63.1 ;
        RECT 36.894 63.098 53.862 63.146 ;
        RECT 36.848 63.144 53.816 63.192 ;
        RECT 36.802 63.19 53.77 63.238 ;
        RECT 36.756 63.236 53.724 63.284 ;
        RECT 36.71 63.282 53.678 63.33 ;
        RECT 36.664 63.328 53.632 63.376 ;
        RECT 36.618 63.374 53.586 63.422 ;
        RECT 36.572 63.42 53.54 63.468 ;
        RECT 36.526 63.466 53.494 63.514 ;
        RECT 36.48 63.512 53.448 63.56 ;
        RECT 36.434 63.558 53.402 63.606 ;
        RECT 36.388 63.604 53.356 63.652 ;
        RECT 36.342 63.65 53.31 63.698 ;
        RECT 36.296 63.696 53.264 63.744 ;
        RECT 36.25 63.742 53.218 63.79 ;
        RECT 36.204 63.788 53.172 63.836 ;
        RECT 36.158 63.834 53.126 63.882 ;
        RECT 36.112 63.88 53.08 63.928 ;
        RECT 36.066 63.926 53.034 63.974 ;
        RECT 36.02 63.972 52.988 64.02 ;
        RECT 35.974 64.018 52.942 64.066 ;
        RECT 35.928 64.064 52.896 64.112 ;
        RECT 35.882 64.11 52.85 64.158 ;
        RECT 35.836 64.156 52.804 64.204 ;
        RECT 35.79 64.202 52.758 64.25 ;
        RECT 35.744 64.248 52.712 64.296 ;
        RECT 35.698 64.294 52.666 64.342 ;
        RECT 35.652 64.34 52.62 64.388 ;
        RECT 35.606 64.386 52.574 64.434 ;
        RECT 35.56 64.432 52.528 64.48 ;
        RECT 35.514 64.478 52.482 64.526 ;
        RECT 35.468 64.524 52.436 64.572 ;
        RECT 35.422 64.57 52.39 64.618 ;
        RECT 35.376 64.616 52.344 64.664 ;
        RECT 35.33 64.662 52.298 64.71 ;
        RECT 35.284 64.708 52.252 64.756 ;
        RECT 35.238 64.754 52.206 64.802 ;
        RECT 35.192 64.8 52.16 64.848 ;
        RECT 35.146 64.846 52.114 64.894 ;
        RECT 35.1 64.892 52.068 64.94 ;
        RECT 35.054 64.938 52.022 64.986 ;
        RECT 35.008 64.984 51.976 65.032 ;
        RECT 34.962 65.03 51.93 65.078 ;
        RECT 34.916 65.076 51.884 65.124 ;
        RECT 34.87 65.122 51.838 65.17 ;
        RECT 34.824 65.168 51.792 65.216 ;
        RECT 34.778 65.214 51.746 65.262 ;
        RECT 34.732 65.26 51.7 65.308 ;
        RECT 34.686 65.306 51.654 65.354 ;
        RECT 34.64 65.352 51.608 65.4 ;
        RECT 34.594 65.398 51.562 65.446 ;
        RECT 34.548 65.444 51.516 65.492 ;
        RECT 34.502 65.49 51.47 65.538 ;
        RECT 34.456 65.536 51.424 65.584 ;
        RECT 34.41 65.582 51.378 65.63 ;
        RECT 34.364 65.628 51.332 65.676 ;
        RECT 34.318 65.674 51.286 65.722 ;
        RECT 34.272 65.72 51.24 65.768 ;
        RECT 34.226 65.766 51.194 65.814 ;
        RECT 34.18 65.812 51.148 65.86 ;
        RECT 34.134 65.858 51.102 65.906 ;
        RECT 34.088 65.904 51.056 65.952 ;
        RECT 34.042 65.95 51.01 65.998 ;
        RECT 33.996 65.996 50.964 66.044 ;
        RECT 33.95 66.042 50.918 66.09 ;
        RECT 33.904 66.088 50.872 66.136 ;
        RECT 33.858 66.134 50.826 66.182 ;
        RECT 33.812 66.18 50.78 66.228 ;
        RECT 33.766 66.226 50.734 66.274 ;
        RECT 33.72 66.272 50.688 66.32 ;
        RECT 33.674 66.318 50.642 66.366 ;
        RECT 33.628 66.364 50.596 66.412 ;
        RECT 33.582 66.41 50.55 66.458 ;
        RECT 33.536 66.456 50.504 66.504 ;
        RECT 33.49 66.502 50.458 66.55 ;
        RECT 33.444 66.548 50.412 66.596 ;
        RECT 33.398 66.594 50.366 66.642 ;
        RECT 33.352 66.64 50.32 66.688 ;
        RECT 33.306 66.686 50.274 66.734 ;
        RECT 33.26 66.732 50.228 66.78 ;
        RECT 33.214 66.778 50.182 66.826 ;
        RECT 33.168 66.824 50.136 66.872 ;
        RECT 33.122 66.87 50.09 66.918 ;
        RECT 33.076 66.916 50.044 66.964 ;
        RECT 33.03 66.962 49.998 67.01 ;
        RECT 32.984 67.008 49.952 67.056 ;
        RECT 32.938 67.054 49.906 67.102 ;
        RECT 32.892 67.1 49.86 67.148 ;
        RECT 32.846 67.146 49.814 67.194 ;
        RECT 32.8 67.192 49.768 67.24 ;
        RECT 32.754 67.238 49.722 67.286 ;
        RECT 32.708 67.284 49.676 67.332 ;
        RECT 32.662 67.33 49.63 67.378 ;
        RECT 32.616 67.376 49.584 67.424 ;
        RECT 32.57 67.422 49.538 67.47 ;
        RECT 32.524 67.468 49.492 67.516 ;
        RECT 32.478 67.514 49.446 67.562 ;
        RECT 32.432 67.56 49.4 67.608 ;
        RECT 32.386 67.606 49.354 67.654 ;
        RECT 32.34 67.652 49.308 67.7 ;
        RECT 32.294 67.698 49.262 67.746 ;
        RECT 32.248 67.744 49.216 67.792 ;
        RECT 32.202 67.79 49.17 67.838 ;
        RECT 32.156 67.836 49.124 67.884 ;
        RECT 32.11 67.882 49.078 67.93 ;
        RECT 32.064 67.928 49.032 67.976 ;
        RECT 32.018 67.974 48.986 68.022 ;
        RECT 31.972 68.02 48.94 68.068 ;
        RECT 31.926 68.066 48.894 68.114 ;
        RECT 31.88 68.112 48.848 68.16 ;
        RECT 31.834 68.158 48.802 68.206 ;
        RECT 31.788 68.204 48.756 68.252 ;
        RECT 31.742 68.25 48.71 68.298 ;
        RECT 31.696 68.296 48.664 68.344 ;
        RECT 31.65 68.342 48.618 68.39 ;
        RECT 31.604 68.388 48.572 68.436 ;
        RECT 31.558 68.434 48.526 68.482 ;
        RECT 31.512 68.48 48.48 68.528 ;
        RECT 31.466 68.526 48.434 68.574 ;
        RECT 31.42 68.572 48.388 68.62 ;
        RECT 31.374 68.618 48.342 68.666 ;
        RECT 31.328 68.664 48.296 68.712 ;
        RECT 31.282 68.71 48.25 68.758 ;
        RECT 31.236 68.756 48.204 68.804 ;
        RECT 31.19 68.802 48.158 68.85 ;
        RECT 31.144 68.848 48.112 68.896 ;
        RECT 31.098 68.894 48.066 68.942 ;
        RECT 31.052 68.94 48.02 68.988 ;
        RECT 31.006 68.986 47.974 69.034 ;
        RECT 30.96 69.032 47.928 69.08 ;
        RECT 30.914 69.078 47.882 69.126 ;
        RECT 30.868 69.124 47.836 69.172 ;
        RECT 30.822 69.17 47.79 69.218 ;
        RECT 30.776 69.216 47.744 69.264 ;
        RECT 30.73 69.262 47.698 69.31 ;
        RECT 30.684 69.308 47.652 69.356 ;
        RECT 30.638 69.354 47.606 69.402 ;
        RECT 30.592 69.4 47.56 69.448 ;
        RECT 30.546 69.446 47.514 69.494 ;
        RECT 30.5 69.492 47.468 69.54 ;
        RECT 30.5 69.492 47.422 69.586 ;
        RECT 30.5 69.492 47.376 69.632 ;
        RECT 30.5 69.492 47.33 69.678 ;
        RECT 30.5 69.492 47.284 69.724 ;
        RECT 30.5 69.492 47.238 69.77 ;
        RECT 30.5 69.492 47.192 69.816 ;
        RECT 30.5 69.492 47.146 69.862 ;
        RECT 30.5 69.492 47.1 69.908 ;
        RECT 30.5 69.492 47.054 69.954 ;
        RECT 30.5 69.492 47.008 70 ;
        RECT 30.5 69.492 46.962 70.046 ;
        RECT 30.5 69.492 46.916 70.092 ;
        RECT 30.5 69.492 46.87 70.138 ;
        RECT 30.5 69.492 46.824 70.184 ;
        RECT 30.5 69.492 46.778 70.23 ;
        RECT 30.5 69.492 46.732 70.276 ;
        RECT 30.5 69.492 46.686 70.322 ;
        RECT 30.5 69.492 46.64 70.368 ;
        RECT 30.5 69.492 46.594 70.414 ;
        RECT 30.5 69.492 46.548 70.46 ;
        RECT 30.5 69.492 46.502 70.506 ;
        RECT 30.5 69.492 46.456 70.552 ;
        RECT 30.5 69.492 46.41 70.598 ;
        RECT 30.5 69.492 46.364 70.644 ;
        RECT 30.5 69.492 46.318 70.69 ;
        RECT 30.5 69.492 46.272 70.736 ;
        RECT 30.5 69.492 46.226 70.782 ;
        RECT 30.5 69.492 46.18 70.828 ;
        RECT 30.5 69.492 46.134 70.874 ;
        RECT 30.5 69.492 46.088 70.92 ;
        RECT 30.5 69.492 46.042 70.966 ;
        RECT 30.5 69.492 45.996 71.012 ;
        RECT 30.5 69.492 45.95 71.058 ;
        RECT 30.5 69.492 45.904 71.104 ;
        RECT 30.5 69.492 45.858 71.15 ;
        RECT 30.5 69.492 45.812 71.196 ;
        RECT 30.5 69.492 45.766 71.242 ;
        RECT 30.5 69.492 45.72 71.288 ;
        RECT 30.5 69.492 45.674 71.334 ;
        RECT 30.5 69.492 45.628 71.38 ;
        RECT 30.5 69.492 45.582 71.426 ;
        RECT 30.5 69.492 45.536 71.472 ;
        RECT 30.5 69.492 45.49 71.518 ;
        RECT 30.5 69.492 45.444 71.564 ;
        RECT 30.5 69.492 45.398 71.61 ;
        RECT 30.5 69.492 45.352 71.656 ;
        RECT 30.5 69.492 45.306 71.702 ;
        RECT 30.5 69.492 45.26 71.748 ;
        RECT 30.5 69.492 45.214 71.794 ;
        RECT 30.5 69.492 45.168 71.84 ;
        RECT 30.5 69.492 45.122 71.886 ;
        RECT 30.5 69.492 45.076 71.932 ;
        RECT 30.5 69.492 45.03 71.978 ;
        RECT 30.5 69.492 44.984 72.024 ;
        RECT 30.5 69.492 44.938 72.07 ;
        RECT 30.5 69.492 44.892 72.116 ;
        RECT 30.5 69.492 44.846 72.162 ;
        RECT 30.5 69.492 44.8 72.208 ;
        RECT 30.5 69.492 44.754 72.254 ;
        RECT 30.5 69.492 44.708 72.3 ;
        RECT 30.5 69.492 44.662 72.346 ;
        RECT 30.5 69.492 44.616 72.392 ;
        RECT 30.5 69.492 44.57 72.438 ;
        RECT 30.5 69.492 44.524 72.484 ;
        RECT 30.5 69.492 44.478 72.53 ;
        RECT 30.5 69.492 44.432 72.576 ;
        RECT 30.5 69.492 44.386 72.622 ;
        RECT 30.5 69.492 44.34 72.668 ;
        RECT 30.5 69.492 44.294 72.714 ;
        RECT 30.5 69.492 44.248 72.76 ;
        RECT 30.5 69.492 44.202 72.806 ;
        RECT 30.5 69.492 44.156 72.852 ;
        RECT 30.5 69.492 44.11 72.898 ;
        RECT 30.5 69.492 44.064 72.944 ;
        RECT 30.5 69.492 44.018 72.99 ;
        RECT 30.5 69.492 43.972 73.036 ;
        RECT 30.5 69.492 43.926 73.082 ;
        RECT 30.5 69.492 43.88 73.128 ;
        RECT 30.5 69.492 43.834 73.174 ;
        RECT 30.5 69.492 43.788 73.22 ;
        RECT 30.5 69.492 43.742 73.266 ;
        RECT 30.5 69.492 43.696 73.312 ;
        RECT 30.5 69.492 43.65 73.358 ;
        RECT 30.5 69.492 43.604 73.404 ;
        RECT 30.5 69.492 43.558 73.45 ;
        RECT 30.5 69.492 43.512 73.496 ;
        RECT 30.5 69.492 43.466 73.542 ;
        RECT 30.5 69.492 43.42 73.588 ;
        RECT 30.5 69.492 43.374 73.634 ;
        RECT 30.5 69.492 43.328 73.68 ;
        RECT 30.5 69.492 43.282 73.726 ;
        RECT 30.5 69.492 43.236 73.772 ;
        RECT 30.5 69.492 43.19 73.818 ;
        RECT 30.5 69.492 43.144 73.864 ;
        RECT 30.5 69.492 43.098 73.91 ;
        RECT 30.5 69.492 43.052 73.956 ;
        RECT 30.5 69.492 43.006 74.002 ;
        RECT 30.5 69.492 42.96 74.048 ;
        RECT 30.5 69.492 42.914 74.094 ;
        RECT 30.5 69.492 42.868 74.14 ;
        RECT 30.5 69.492 42.822 74.186 ;
        RECT 30.5 69.492 42.776 74.232 ;
        RECT 30.5 69.492 42.73 74.278 ;
        RECT 30.5 69.492 42.684 74.324 ;
        RECT 30.5 69.492 42.638 74.37 ;
        RECT 30.5 69.492 42.592 74.416 ;
        RECT 30.5 69.492 42.546 74.462 ;
        RECT 30.5 69.492 42.5 110 ;
        RECT 76.265 44 110 56 ;
        RECT 59.312 60.93 76.265 60.983 ;
        RECT 59.358 60.884 76.311 60.947 ;
        RECT 76.24 44.012 76.265 60.983 ;
        RECT 59.404 60.838 76.357 60.901 ;
        RECT 76.194 44.048 76.24 61.018 ;
        RECT 59.266 60.976 76.194 61.064 ;
        RECT 59.45 60.792 76.403 60.855 ;
        RECT 76.148 44.094 76.194 61.064 ;
        RECT 59.22 61.022 76.148 61.11 ;
        RECT 59.496 60.746 76.449 60.809 ;
        RECT 76.102 44.14 76.148 61.11 ;
        RECT 59.174 61.068 76.102 61.156 ;
        RECT 59.542 60.7 76.495 60.763 ;
        RECT 76.056 44.186 76.102 61.156 ;
        RECT 59.128 61.114 76.056 61.202 ;
        RECT 59.588 60.654 76.541 60.717 ;
        RECT 76.01 44.232 76.056 61.202 ;
        RECT 59.082 61.16 76.01 61.248 ;
        RECT 59.634 60.608 76.587 60.671 ;
        RECT 75.964 44.278 76.01 61.248 ;
        RECT 59.036 61.206 75.964 61.294 ;
        RECT 59.68 60.562 76.633 60.625 ;
        RECT 75.918 44.324 75.964 61.294 ;
        RECT 58.99 61.252 75.918 61.34 ;
        RECT 59.726 60.516 76.679 60.579 ;
        RECT 75.872 44.37 75.918 61.34 ;
        RECT 58.944 61.298 75.872 61.386 ;
        RECT 59.772 60.47 76.725 60.533 ;
        RECT 75.826 44.416 75.872 61.386 ;
        RECT 58.898 61.344 75.826 61.432 ;
        RECT 59.818 60.424 76.771 60.487 ;
        RECT 75.78 44.462 75.826 61.432 ;
        RECT 58.852 61.39 75.78 61.478 ;
        RECT 59.864 60.378 76.817 60.441 ;
        RECT 75.734 44.508 75.78 61.478 ;
        RECT 58.806 61.436 75.734 61.524 ;
        RECT 59.91 60.332 76.863 60.395 ;
        RECT 75.688 44.554 75.734 61.524 ;
        RECT 58.76 61.482 75.688 61.57 ;
        RECT 59.956 60.286 76.909 60.349 ;
      LAYER MET3 ;
        RECT 70.814 69.423 79.278 69.485 ;
        RECT 77.852 62.385 110 63.5 ;
        RECT 79.232 61.005 79.278 69.485 ;
        RECT 70.768 69.469 79.232 69.531 ;
        RECT 77.898 62.339 110 63.5 ;
        RECT 79.186 61.051 79.232 69.531 ;
        RECT 70.722 69.515 79.186 69.577 ;
        RECT 77.944 62.293 110 63.5 ;
        RECT 79.14 61.097 79.186 69.577 ;
        RECT 70.676 69.561 79.14 69.623 ;
        RECT 77.99 62.247 110 63.5 ;
        RECT 79.094 61.143 79.14 69.623 ;
        RECT 70.63 69.607 79.094 69.669 ;
        RECT 78.036 62.201 110 63.5 ;
        RECT 79.048 61.189 79.094 69.669 ;
        RECT 70.584 69.653 79.048 69.715 ;
        RECT 78.082 62.155 110 63.5 ;
        RECT 79.002 61.235 79.048 69.715 ;
        RECT 70.538 69.699 79.002 69.761 ;
        RECT 78.128 62.109 110 63.5 ;
        RECT 78.956 61.281 79.002 69.761 ;
        RECT 70.492 69.745 78.956 69.807 ;
        RECT 78.174 62.063 110 63.5 ;
        RECT 78.91 61.327 78.956 69.807 ;
        RECT 70.446 69.791 78.91 69.853 ;
        RECT 78.22 62.017 110 63.5 ;
        RECT 78.864 61.373 78.91 69.853 ;
        RECT 70.4 69.837 78.864 69.899 ;
        RECT 78.266 61.971 110 63.5 ;
        RECT 78.818 61.419 78.864 69.899 ;
        RECT 70.354 69.883 78.818 69.945 ;
        RECT 78.312 61.925 110 63.5 ;
        RECT 78.772 61.465 78.818 69.945 ;
        RECT 70.308 69.929 78.772 69.991 ;
        RECT 78.358 61.879 110 63.5 ;
        RECT 78.726 61.511 78.772 69.991 ;
        RECT 70.262 69.975 78.726 70.037 ;
        RECT 78.404 61.833 110 63.5 ;
        RECT 78.68 61.557 78.726 70.037 ;
        RECT 70.216 70.021 78.68 70.083 ;
        RECT 78.45 61.787 110 63.5 ;
        RECT 78.634 61.603 78.68 70.083 ;
        RECT 70.17 70.067 78.634 70.129 ;
        RECT 78.496 61.741 110 63.5 ;
        RECT 78.588 61.649 78.634 70.129 ;
        RECT 70.124 70.113 78.588 70.175 ;
        RECT 78.542 61.695 110 63.5 ;
        RECT 70.078 70.159 78.542 70.221 ;
        RECT 70.032 70.205 78.496 70.267 ;
        RECT 69.986 70.251 78.45 70.313 ;
        RECT 69.94 70.297 78.404 70.359 ;
        RECT 69.894 70.343 78.358 70.405 ;
        RECT 69.848 70.389 78.312 70.451 ;
        RECT 69.802 70.435 78.266 70.497 ;
        RECT 69.756 70.481 78.22 70.543 ;
        RECT 69.71 70.527 78.174 70.589 ;
        RECT 69.664 70.573 78.128 70.635 ;
        RECT 69.618 70.619 78.082 70.681 ;
        RECT 69.572 70.665 78.036 70.727 ;
        RECT 69.526 70.711 77.99 70.773 ;
        RECT 69.48 70.757 77.944 70.819 ;
        RECT 69.434 70.803 77.898 70.865 ;
        RECT 69.388 70.849 77.852 70.911 ;
        RECT 69.342 70.895 77.806 70.957 ;
        RECT 69.296 70.941 77.76 71.003 ;
        RECT 69.25 70.987 77.714 71.049 ;
        RECT 69.204 71.033 77.668 71.095 ;
        RECT 69.158 71.079 77.622 71.141 ;
        RECT 69.112 71.125 77.576 71.187 ;
        RECT 69.066 71.171 77.53 71.233 ;
        RECT 69.02 71.217 77.484 71.279 ;
        RECT 68.974 71.263 77.438 71.325 ;
        RECT 68.928 71.309 77.392 71.371 ;
        RECT 68.882 71.355 77.346 71.417 ;
        RECT 68.836 71.401 77.3 71.463 ;
        RECT 68.79 71.447 77.254 71.509 ;
        RECT 68.744 71.493 77.208 71.555 ;
        RECT 68.698 71.539 77.162 71.601 ;
        RECT 68.652 71.585 77.116 71.647 ;
        RECT 68.606 71.631 77.07 71.693 ;
        RECT 68.56 71.677 77.024 71.739 ;
        RECT 68.514 71.723 76.978 71.785 ;
        RECT 68.468 71.769 76.932 71.831 ;
        RECT 68.422 71.815 76.886 71.877 ;
        RECT 68.376 71.861 76.84 71.923 ;
        RECT 68.33 71.907 76.794 71.969 ;
        RECT 68.284 71.953 76.748 72.015 ;
        RECT 68.238 71.999 76.702 72.061 ;
        RECT 68.192 72.045 76.656 72.107 ;
        RECT 68.146 72.091 76.61 72.153 ;
        RECT 68.1 72.137 76.564 72.199 ;
        RECT 68.054 72.183 76.518 72.245 ;
        RECT 68.008 72.229 76.472 72.291 ;
        RECT 67.962 72.275 76.426 72.337 ;
        RECT 67.916 72.321 76.38 72.383 ;
        RECT 67.87 72.367 76.334 72.429 ;
        RECT 67.824 72.413 76.288 72.475 ;
        RECT 67.778 72.459 76.242 72.521 ;
        RECT 67.732 72.505 76.196 72.567 ;
        RECT 67.686 72.551 76.15 72.613 ;
        RECT 67.64 72.597 76.104 72.659 ;
        RECT 67.594 72.643 76.058 72.705 ;
        RECT 67.548 72.689 76.012 72.751 ;
        RECT 67.502 72.735 75.966 72.797 ;
        RECT 67.456 72.781 75.92 72.843 ;
        RECT 67.41 72.827 75.874 72.889 ;
        RECT 67.364 72.873 75.828 72.935 ;
        RECT 67.318 72.919 75.782 72.981 ;
        RECT 67.272 72.965 75.736 73.027 ;
        RECT 67.226 73.011 75.69 73.073 ;
        RECT 67.18 73.057 75.644 73.119 ;
        RECT 67.134 73.103 75.598 73.165 ;
        RECT 67.088 73.149 75.552 73.211 ;
        RECT 67.042 73.195 75.506 73.257 ;
        RECT 66.996 73.241 75.46 73.303 ;
        RECT 66.95 73.287 75.414 73.349 ;
        RECT 66.904 73.333 75.368 73.395 ;
        RECT 66.858 73.379 75.322 73.441 ;
        RECT 66.812 73.425 75.276 73.487 ;
        RECT 66.766 73.471 75.23 73.533 ;
        RECT 66.72 73.517 75.184 73.579 ;
        RECT 66.674 73.563 75.138 73.625 ;
        RECT 66.628 73.609 75.092 73.671 ;
        RECT 66.582 73.655 75.046 73.717 ;
        RECT 66.536 73.701 75 73.763 ;
        RECT 66.49 73.747 74.954 73.809 ;
        RECT 66.444 73.793 74.908 73.855 ;
        RECT 66.398 73.839 74.862 73.901 ;
        RECT 66.352 73.885 74.816 73.947 ;
        RECT 66.306 73.931 74.77 73.993 ;
        RECT 66.26 73.977 74.724 74.039 ;
        RECT 66.214 74.023 74.678 74.085 ;
        RECT 66.168 74.069 74.632 74.131 ;
        RECT 66.122 74.115 74.586 74.177 ;
        RECT 66.076 74.161 74.54 74.223 ;
        RECT 66.03 74.207 74.494 74.269 ;
        RECT 65.984 74.253 74.448 74.315 ;
        RECT 65.938 74.299 74.402 74.361 ;
        RECT 65.892 74.345 74.356 74.407 ;
        RECT 65.846 74.391 74.31 74.453 ;
        RECT 65.8 74.437 74.264 74.499 ;
        RECT 65.754 74.483 74.218 74.545 ;
        RECT 65.708 74.529 74.172 74.591 ;
        RECT 65.662 74.575 74.126 74.637 ;
        RECT 65.616 74.621 74.08 74.683 ;
        RECT 65.57 74.667 74.034 74.729 ;
        RECT 65.524 74.713 73.988 74.775 ;
        RECT 65.478 74.759 73.942 74.821 ;
        RECT 65.432 74.805 73.896 74.867 ;
        RECT 65.386 74.851 73.85 74.913 ;
        RECT 65.34 74.897 73.804 74.959 ;
        RECT 65.294 74.943 73.758 75.005 ;
        RECT 65.248 74.989 73.712 75.051 ;
        RECT 65.202 75.035 73.666 75.097 ;
        RECT 65.156 75.081 73.62 75.143 ;
        RECT 65.11 75.127 73.574 75.189 ;
        RECT 65.064 75.173 73.528 75.235 ;
        RECT 65.018 75.219 73.482 75.281 ;
        RECT 64.972 75.265 73.436 75.327 ;
        RECT 64.926 75.311 73.39 75.373 ;
        RECT 64.88 75.357 73.344 75.419 ;
        RECT 64.834 75.403 73.298 75.465 ;
        RECT 64.788 75.449 73.252 75.511 ;
        RECT 64.742 75.495 73.206 75.557 ;
        RECT 64.696 75.541 73.16 75.603 ;
        RECT 64.65 75.587 73.114 75.649 ;
        RECT 64.604 75.633 73.068 75.695 ;
        RECT 64.558 75.679 73.022 75.741 ;
        RECT 64.512 75.725 72.976 75.787 ;
        RECT 64.466 75.771 72.93 75.833 ;
        RECT 64.42 75.817 72.884 75.879 ;
        RECT 64.374 75.863 72.838 75.925 ;
        RECT 64.328 75.909 72.792 75.971 ;
        RECT 64.282 75.955 72.746 76.017 ;
        RECT 64.236 76.001 72.7 76.063 ;
        RECT 64.19 76.047 72.654 76.109 ;
        RECT 64.144 76.093 72.608 76.155 ;
        RECT 64.098 76.139 72.562 76.201 ;
        RECT 64.052 76.185 72.516 76.247 ;
        RECT 64.006 76.231 72.47 76.293 ;
        RECT 63.96 76.277 72.424 76.339 ;
        RECT 63.914 76.323 72.378 76.385 ;
        RECT 63.868 76.369 72.332 76.431 ;
        RECT 63.822 76.415 72.286 76.477 ;
        RECT 63.776 76.461 72.24 76.523 ;
        RECT 63.73 76.507 72.194 76.569 ;
        RECT 63.684 76.553 72.148 76.615 ;
        RECT 63.638 76.599 72.102 76.661 ;
        RECT 63.592 76.645 72.056 76.707 ;
        RECT 63.546 76.691 72.01 76.753 ;
        RECT 63.5 76.737 71.964 76.799 ;
        RECT 63.48 76.77 71.918 76.845 ;
        RECT 63.434 76.803 71.872 76.891 ;
        RECT 63.388 76.849 71.826 76.937 ;
        RECT 63.342 76.895 71.78 76.983 ;
        RECT 63.296 76.941 71.734 77.029 ;
        RECT 63.25 76.987 71.688 77.075 ;
        RECT 63.204 77.033 71.642 77.121 ;
        RECT 63.158 77.079 71.596 77.167 ;
        RECT 63.112 77.125 71.55 77.213 ;
        RECT 63.066 77.171 71.504 77.259 ;
        RECT 63.02 77.217 71.458 77.305 ;
        RECT 62.974 77.263 71.412 77.351 ;
        RECT 62.928 77.309 71.366 77.397 ;
        RECT 62.882 77.355 71.32 77.443 ;
        RECT 62.836 77.401 71.274 77.489 ;
        RECT 62.79 77.447 71.228 77.535 ;
        RECT 62.744 77.493 71.182 77.581 ;
        RECT 62.698 77.539 71.136 77.627 ;
        RECT 62.652 77.585 71.09 77.673 ;
        RECT 62.606 77.631 71.044 77.719 ;
        RECT 62.56 77.677 70.998 77.765 ;
        RECT 62.514 77.723 70.952 77.811 ;
        RECT 62.468 77.769 70.906 77.857 ;
        RECT 62.422 77.815 70.86 77.903 ;
        RECT 62.376 77.861 70.814 77.949 ;
        RECT 62.33 77.907 70.768 77.995 ;
        RECT 62.284 77.953 70.722 78.041 ;
        RECT 62.238 77.999 70.676 78.087 ;
        RECT 62.192 78.045 70.63 78.133 ;
        RECT 62.146 78.091 70.584 78.179 ;
        RECT 62.1 78.137 70.538 78.225 ;
        RECT 62.054 78.183 70.492 78.271 ;
        RECT 62.008 78.229 70.446 78.317 ;
        RECT 61.962 78.275 70.4 78.363 ;
        RECT 61.916 78.321 70.354 78.409 ;
        RECT 61.87 78.367 70.308 78.455 ;
        RECT 61.824 78.413 70.262 78.501 ;
        RECT 61.778 78.459 70.216 78.547 ;
        RECT 61.732 78.505 70.17 78.593 ;
        RECT 61.686 78.551 70.124 78.639 ;
        RECT 61.64 78.597 70.078 78.685 ;
        RECT 61.594 78.643 70.032 78.731 ;
        RECT 61.548 78.689 69.986 78.777 ;
        RECT 61.502 78.735 69.94 78.823 ;
        RECT 61.456 78.781 69.894 78.869 ;
        RECT 61.41 78.827 69.848 78.915 ;
        RECT 61.364 78.873 69.802 78.961 ;
        RECT 61.318 78.919 69.756 79.007 ;
        RECT 61.272 78.965 69.71 79.053 ;
        RECT 61.226 79.011 69.664 79.099 ;
        RECT 61.18 79.057 69.618 79.145 ;
        RECT 61.134 79.103 69.572 79.191 ;
        RECT 61.088 79.149 69.526 79.237 ;
        RECT 61.042 79.195 69.48 79.283 ;
        RECT 60.996 79.241 69.434 79.329 ;
        RECT 60.95 79.287 69.388 79.375 ;
        RECT 60.904 79.333 69.342 79.421 ;
        RECT 60.858 79.379 69.296 79.467 ;
        RECT 60.812 79.425 69.25 79.513 ;
        RECT 60.766 79.471 69.204 79.559 ;
        RECT 60.72 79.517 69.158 79.605 ;
        RECT 60.674 79.563 69.112 79.651 ;
        RECT 60.628 79.609 69.066 79.697 ;
        RECT 60.582 79.655 69.02 79.743 ;
        RECT 60.536 79.701 68.974 79.789 ;
        RECT 60.49 79.747 68.928 79.835 ;
        RECT 60.444 79.793 68.882 79.881 ;
        RECT 60.398 79.839 68.836 79.927 ;
        RECT 60.352 79.885 68.79 79.973 ;
        RECT 60.306 79.931 68.744 80.019 ;
        RECT 60.26 79.977 68.698 80.065 ;
        RECT 60.214 80.023 68.652 80.111 ;
        RECT 60.168 80.069 68.606 80.157 ;
        RECT 60.122 80.115 68.56 80.203 ;
        RECT 60.076 80.161 68.514 80.249 ;
        RECT 60.03 80.207 68.468 80.295 ;
        RECT 59.984 80.253 68.422 80.341 ;
        RECT 59.938 80.299 68.376 80.387 ;
        RECT 59.892 80.345 68.33 80.433 ;
        RECT 59.846 80.391 68.284 80.479 ;
        RECT 59.8 80.437 68.238 80.525 ;
        RECT 59.754 80.483 68.192 80.571 ;
        RECT 59.708 80.529 68.146 80.617 ;
        RECT 59.662 80.575 68.1 80.663 ;
        RECT 59.616 80.621 68.054 80.709 ;
        RECT 59.57 80.667 68.008 80.755 ;
        RECT 59.524 80.713 67.962 80.801 ;
        RECT 59.478 80.759 67.916 80.847 ;
        RECT 59.432 80.805 67.87 80.893 ;
        RECT 59.386 80.851 67.824 80.939 ;
        RECT 59.34 80.897 67.778 80.985 ;
        RECT 59.294 80.943 67.732 81.031 ;
        RECT 59.248 80.989 67.686 81.077 ;
        RECT 59.202 81.035 67.64 81.123 ;
        RECT 59.156 81.081 67.594 81.169 ;
        RECT 59.11 81.127 67.548 81.215 ;
        RECT 59.064 81.173 67.502 81.261 ;
        RECT 59.018 81.219 67.456 81.307 ;
        RECT 58.972 81.265 67.41 81.353 ;
        RECT 58.926 81.311 67.364 81.399 ;
        RECT 58.88 81.357 67.318 81.445 ;
        RECT 58.834 81.403 67.272 81.491 ;
        RECT 58.788 81.449 67.226 81.537 ;
        RECT 58.742 81.495 67.18 81.583 ;
        RECT 58.696 81.541 67.134 81.629 ;
        RECT 58.65 81.587 67.088 81.675 ;
        RECT 58.604 81.633 67.042 81.721 ;
        RECT 58.558 81.679 66.996 81.767 ;
        RECT 58.512 81.725 66.95 81.813 ;
        RECT 58.466 81.771 66.904 81.859 ;
        RECT 58.42 81.817 66.858 81.905 ;
        RECT 58.374 81.863 66.812 81.951 ;
        RECT 58.328 81.909 66.766 81.997 ;
        RECT 58.282 81.955 66.72 82.043 ;
        RECT 58.236 82.001 66.674 82.089 ;
        RECT 58.19 82.047 66.628 82.135 ;
        RECT 58.144 82.093 66.582 82.181 ;
        RECT 58.098 82.139 66.536 82.227 ;
        RECT 58.052 82.185 66.49 82.273 ;
        RECT 58.006 82.231 66.444 82.319 ;
        RECT 57.96 82.277 66.398 82.365 ;
        RECT 57.914 82.323 66.352 82.411 ;
        RECT 57.868 82.369 66.306 82.457 ;
        RECT 57.822 82.415 66.26 82.503 ;
        RECT 57.776 82.461 66.214 82.549 ;
        RECT 57.73 82.507 66.168 82.595 ;
        RECT 57.684 82.553 66.122 82.641 ;
        RECT 57.638 82.599 66.076 82.687 ;
        RECT 57.592 82.645 66.03 82.733 ;
        RECT 57.546 82.691 65.984 82.779 ;
        RECT 57.5 82.737 65.938 82.825 ;
        RECT 57.5 82.737 65.892 82.871 ;
        RECT 57.5 82.737 65.846 82.917 ;
        RECT 57.5 82.737 65.8 82.963 ;
        RECT 57.5 82.737 65.754 83.009 ;
        RECT 57.5 82.737 65.708 83.055 ;
        RECT 57.5 82.737 65.662 83.101 ;
        RECT 57.5 82.737 65.616 83.147 ;
        RECT 57.5 82.737 65.57 83.193 ;
        RECT 57.5 82.737 65.524 83.239 ;
        RECT 57.5 82.737 65.478 83.285 ;
        RECT 57.5 82.737 65.432 83.331 ;
        RECT 57.5 82.737 65.386 83.377 ;
        RECT 57.5 82.737 65.34 83.423 ;
        RECT 57.5 82.737 65.294 83.469 ;
        RECT 57.5 82.737 65.248 83.515 ;
        RECT 57.5 82.737 65.202 83.561 ;
        RECT 57.5 82.737 65.156 83.607 ;
        RECT 57.5 82.737 65.11 83.653 ;
        RECT 57.5 82.737 65.064 83.699 ;
        RECT 57.5 82.737 65.018 83.745 ;
        RECT 57.5 82.737 64.972 83.791 ;
        RECT 57.5 82.737 64.926 83.837 ;
        RECT 57.5 82.737 64.88 83.883 ;
        RECT 57.5 82.737 64.834 83.929 ;
        RECT 57.5 82.737 64.788 83.975 ;
        RECT 57.5 82.737 64.742 84.021 ;
        RECT 57.5 82.737 64.696 84.067 ;
        RECT 57.5 82.737 64.65 84.113 ;
        RECT 57.5 82.737 64.604 84.159 ;
        RECT 57.5 82.737 64.558 84.205 ;
        RECT 57.5 82.737 64.512 84.251 ;
        RECT 57.5 82.737 64.466 84.297 ;
        RECT 57.5 82.737 64.42 84.343 ;
        RECT 57.5 82.737 64.374 84.389 ;
        RECT 57.5 82.737 64.328 84.435 ;
        RECT 57.5 82.737 64.282 84.481 ;
        RECT 57.5 82.737 64.236 84.527 ;
        RECT 57.5 82.737 64.19 84.573 ;
        RECT 57.5 82.737 64.144 84.619 ;
        RECT 57.5 82.737 64.098 84.665 ;
        RECT 57.5 82.737 64.052 84.711 ;
        RECT 57.5 82.737 64.006 84.757 ;
        RECT 57.5 82.737 63.96 84.803 ;
        RECT 57.5 82.737 63.914 84.849 ;
        RECT 57.5 82.737 63.868 84.895 ;
        RECT 57.5 82.737 63.822 84.941 ;
        RECT 57.5 82.737 63.776 84.987 ;
        RECT 57.5 82.737 63.73 85.033 ;
        RECT 57.5 82.737 63.684 85.079 ;
        RECT 57.5 82.737 63.638 85.125 ;
        RECT 57.5 82.737 63.592 85.171 ;
        RECT 57.5 82.737 63.546 85.217 ;
        RECT 57.5 82.737 63.5 110 ;
        RECT 88.365 68.5 110 77 ;
        RECT 79.852 76.99 91.885 77.012 ;
        RECT 76.366 80.476 88.365 80.522 ;
        RECT 76.412 80.43 88.411 80.497 ;
        RECT 88.362 68.501 88.365 80.522 ;
        RECT 76.458 80.384 88.457 80.451 ;
        RECT 88.316 68.526 88.362 80.546 ;
        RECT 76.32 80.522 88.316 80.592 ;
        RECT 76.504 80.338 88.503 80.405 ;
        RECT 88.27 68.572 88.316 80.592 ;
        RECT 76.274 80.568 88.27 80.638 ;
        RECT 76.55 80.292 88.549 80.359 ;
        RECT 88.224 68.618 88.27 80.638 ;
        RECT 76.228 80.614 88.224 80.684 ;
        RECT 76.596 80.246 88.595 80.313 ;
        RECT 88.178 68.664 88.224 80.684 ;
        RECT 76.182 80.66 88.178 80.73 ;
        RECT 76.642 80.2 88.641 80.267 ;
        RECT 88.132 68.71 88.178 80.73 ;
        RECT 76.136 80.706 88.132 80.776 ;
        RECT 76.688 80.154 88.687 80.221 ;
        RECT 88.086 68.756 88.132 80.776 ;
        RECT 76.09 80.752 88.086 80.822 ;
        RECT 76.734 80.108 88.733 80.175 ;
        RECT 88.04 68.802 88.086 80.822 ;
        RECT 76.044 80.798 88.04 80.868 ;
        RECT 76.78 80.062 88.779 80.129 ;
        RECT 87.994 68.848 88.04 80.868 ;
        RECT 75.998 80.844 87.994 80.914 ;
        RECT 76.826 80.016 88.825 80.083 ;
        RECT 87.948 68.894 87.994 80.914 ;
        RECT 75.952 80.89 87.948 80.96 ;
        RECT 76.872 79.97 88.871 80.037 ;
        RECT 87.902 68.94 87.948 80.96 ;
        RECT 75.906 80.936 87.902 81.006 ;
        RECT 76.918 79.924 88.917 79.991 ;
        RECT 87.856 68.986 87.902 81.006 ;
        RECT 75.86 80.982 87.856 81.052 ;
        RECT 76.964 79.883 88.963 79.945 ;
        RECT 87.81 69.032 87.856 81.052 ;
        RECT 75.814 81.028 87.81 81.098 ;
        RECT 77 79.842 89.009 79.899 ;
        RECT 87.764 69.078 87.81 81.098 ;
        RECT 75.768 81.074 87.764 81.144 ;
        RECT 77.046 79.796 89.055 79.853 ;
        RECT 87.718 69.124 87.764 81.144 ;
        RECT 75.722 81.12 87.718 81.19 ;
        RECT 77.092 79.75 89.101 79.807 ;
        RECT 87.672 69.17 87.718 81.19 ;
        RECT 75.676 81.166 87.672 81.236 ;
        RECT 77.138 79.704 89.147 79.761 ;
        RECT 87.626 69.216 87.672 81.236 ;
        RECT 75.63 81.212 87.626 81.282 ;
        RECT 77.184 79.658 89.193 79.715 ;
        RECT 87.58 69.262 87.626 81.282 ;
        RECT 75.584 81.258 87.58 81.328 ;
        RECT 77.23 79.612 89.239 79.669 ;
        RECT 87.534 69.308 87.58 81.328 ;
        RECT 75.538 81.304 87.534 81.374 ;
        RECT 77.276 79.566 89.285 79.623 ;
        RECT 87.488 69.354 87.534 81.374 ;
        RECT 75.492 81.35 87.488 81.42 ;
        RECT 77.322 79.52 89.331 79.577 ;
        RECT 87.442 69.4 87.488 81.42 ;
        RECT 75.446 81.396 87.442 81.466 ;
        RECT 77.368 79.474 89.377 79.531 ;
        RECT 87.396 69.446 87.442 81.466 ;
        RECT 75.4 81.442 87.396 81.512 ;
        RECT 77.414 79.428 89.423 79.485 ;
        RECT 87.35 69.492 87.396 81.512 ;
        RECT 75.354 81.488 87.35 81.558 ;
        RECT 77.46 79.382 89.469 79.439 ;
        RECT 87.304 69.538 87.35 81.558 ;
        RECT 75.308 81.534 87.304 81.604 ;
        RECT 77.506 79.336 89.515 79.393 ;
        RECT 87.258 69.584 87.304 81.604 ;
        RECT 75.262 81.58 87.258 81.65 ;
        RECT 77.552 79.29 89.561 79.347 ;
        RECT 87.212 69.63 87.258 81.65 ;
        RECT 75.216 81.626 87.212 81.696 ;
        RECT 77.598 79.244 89.607 79.301 ;
        RECT 87.166 69.676 87.212 81.696 ;
        RECT 75.17 81.672 87.166 81.742 ;
        RECT 77.644 79.198 89.653 79.255 ;
        RECT 87.12 69.722 87.166 81.742 ;
        RECT 75.124 81.718 87.12 81.788 ;
        RECT 77.69 79.152 89.699 79.209 ;
        RECT 87.074 69.768 87.12 81.788 ;
        RECT 75.078 81.764 87.074 81.834 ;
        RECT 77.736 79.106 89.745 79.163 ;
        RECT 87.028 69.814 87.074 81.834 ;
        RECT 75.032 81.81 87.028 81.88 ;
        RECT 77.782 79.06 89.791 79.117 ;
        RECT 86.982 69.86 87.028 81.88 ;
        RECT 74.986 81.856 86.982 81.926 ;
        RECT 77.828 79.014 89.837 79.071 ;
        RECT 86.936 69.906 86.982 81.926 ;
        RECT 74.94 81.902 86.936 81.972 ;
        RECT 77.874 78.968 89.883 79.025 ;
        RECT 86.89 69.952 86.936 81.972 ;
        RECT 74.894 81.948 86.89 82.018 ;
        RECT 77.92 78.922 89.929 78.979 ;
        RECT 86.844 69.998 86.89 82.018 ;
        RECT 74.848 81.994 86.844 82.064 ;
        RECT 77.966 78.876 89.975 78.933 ;
        RECT 86.798 70.044 86.844 82.064 ;
        RECT 74.802 82.04 86.798 82.11 ;
        RECT 78.012 78.83 90.021 78.887 ;
        RECT 86.752 70.09 86.798 82.11 ;
        RECT 74.756 82.086 86.752 82.156 ;
        RECT 78.058 78.784 90.067 78.841 ;
        RECT 86.706 70.136 86.752 82.156 ;
        RECT 74.71 82.132 86.706 82.202 ;
        RECT 78.104 78.738 90.113 78.795 ;
        RECT 86.66 70.182 86.706 82.202 ;
        RECT 74.664 82.178 86.66 82.248 ;
        RECT 78.15 78.692 90.159 78.749 ;
        RECT 86.614 70.228 86.66 82.248 ;
        RECT 74.618 82.224 86.614 82.294 ;
        RECT 78.196 78.646 90.205 78.703 ;
        RECT 86.568 70.274 86.614 82.294 ;
        RECT 74.572 82.27 86.568 82.34 ;
        RECT 78.242 78.6 90.251 78.657 ;
        RECT 86.522 70.32 86.568 82.34 ;
        RECT 74.526 82.316 86.522 82.386 ;
        RECT 78.288 78.554 90.297 78.611 ;
        RECT 86.476 70.366 86.522 82.386 ;
        RECT 74.48 82.362 86.476 82.432 ;
        RECT 78.334 78.508 90.343 78.565 ;
        RECT 86.43 70.412 86.476 82.432 ;
        RECT 74.434 82.408 86.43 82.478 ;
        RECT 78.38 78.462 90.389 78.519 ;
        RECT 86.384 70.458 86.43 82.478 ;
        RECT 74.388 82.454 86.384 82.524 ;
        RECT 78.426 78.416 90.435 78.473 ;
        RECT 86.338 70.504 86.384 82.524 ;
        RECT 74.342 82.5 86.338 82.57 ;
        RECT 78.472 78.37 90.481 78.427 ;
        RECT 86.292 70.55 86.338 82.57 ;
        RECT 74.296 82.546 86.292 82.616 ;
        RECT 78.518 78.324 90.527 78.381 ;
        RECT 86.246 70.596 86.292 82.616 ;
        RECT 74.25 82.592 86.246 82.662 ;
        RECT 78.564 78.278 90.573 78.335 ;
        RECT 86.2 70.642 86.246 82.662 ;
        RECT 74.204 82.638 86.2 82.708 ;
        RECT 78.61 78.232 90.619 78.289 ;
        RECT 86.154 70.688 86.2 82.708 ;
        RECT 74.158 82.684 86.154 82.754 ;
        RECT 78.656 78.186 90.665 78.243 ;
        RECT 86.108 70.734 86.154 82.754 ;
        RECT 74.112 82.73 86.108 82.8 ;
        RECT 78.702 78.14 90.711 78.197 ;
        RECT 86.062 70.78 86.108 82.8 ;
        RECT 74.066 82.776 86.062 82.846 ;
        RECT 78.748 78.094 90.757 78.151 ;
        RECT 86.016 70.826 86.062 82.846 ;
        RECT 74.02 82.822 86.016 82.892 ;
        RECT 78.794 78.048 90.803 78.105 ;
        RECT 85.97 70.872 86.016 82.892 ;
        RECT 73.974 82.868 85.97 82.938 ;
        RECT 78.84 78.002 90.849 78.059 ;
        RECT 85.924 70.918 85.97 82.938 ;
        RECT 73.928 82.914 85.924 82.984 ;
        RECT 78.886 77.956 90.895 78.013 ;
        RECT 85.878 70.964 85.924 82.984 ;
        RECT 73.882 82.96 85.878 83.03 ;
        RECT 78.932 77.91 90.941 77.967 ;
        RECT 85.832 71.01 85.878 83.03 ;
        RECT 73.836 83.006 85.832 83.076 ;
        RECT 78.978 77.864 90.987 77.921 ;
        RECT 85.786 71.056 85.832 83.076 ;
        RECT 73.79 83.052 85.786 83.122 ;
        RECT 79.024 77.818 91.033 77.875 ;
        RECT 85.74 71.102 85.786 83.122 ;
        RECT 73.744 83.098 85.74 83.168 ;
        RECT 79.07 77.772 91.079 77.829 ;
        RECT 85.694 71.148 85.74 83.168 ;
        RECT 73.698 83.144 85.694 83.214 ;
        RECT 79.116 77.726 91.125 77.783 ;
        RECT 85.648 71.194 85.694 83.214 ;
        RECT 73.652 83.19 85.648 83.26 ;
        RECT 79.162 77.68 91.171 77.737 ;
        RECT 85.602 71.24 85.648 83.26 ;
        RECT 73.606 83.236 85.602 83.306 ;
        RECT 79.208 77.634 91.217 77.691 ;
        RECT 85.556 71.286 85.602 83.306 ;
        RECT 73.56 83.282 85.556 83.352 ;
        RECT 79.254 77.588 91.263 77.645 ;
        RECT 85.51 71.332 85.556 83.352 ;
        RECT 73.514 83.328 85.51 83.398 ;
        RECT 79.3 77.542 91.309 77.599 ;
        RECT 85.464 71.378 85.51 83.398 ;
        RECT 73.468 83.374 85.464 83.444 ;
        RECT 79.346 77.496 91.355 77.553 ;
        RECT 85.418 71.424 85.464 83.444 ;
        RECT 73.422 83.42 85.418 83.49 ;
        RECT 79.392 77.45 91.401 77.507 ;
        RECT 85.372 71.47 85.418 83.49 ;
        RECT 73.376 83.466 85.372 83.536 ;
        RECT 79.438 77.404 91.447 77.461 ;
        RECT 85.326 71.516 85.372 83.536 ;
        RECT 73.33 83.512 85.326 83.582 ;
        RECT 79.484 77.358 91.493 77.415 ;
        RECT 85.28 71.562 85.326 83.582 ;
        RECT 73.284 83.558 85.28 83.628 ;
        RECT 79.53 77.312 91.539 77.369 ;
        RECT 85.234 71.608 85.28 83.628 ;
        RECT 73.238 83.604 85.234 83.674 ;
        RECT 79.576 77.266 91.585 77.323 ;
        RECT 85.188 71.654 85.234 83.674 ;
        RECT 73.192 83.65 85.188 83.72 ;
        RECT 79.622 77.22 91.631 77.277 ;
        RECT 85.142 71.7 85.188 83.72 ;
        RECT 73.146 83.696 85.142 83.766 ;
        RECT 79.668 77.174 91.677 77.231 ;
        RECT 85.096 71.746 85.142 83.766 ;
        RECT 73.1 83.742 85.096 83.812 ;
        RECT 79.714 77.128 91.723 77.185 ;
        RECT 85.05 71.792 85.096 83.812 ;
        RECT 73.054 83.788 85.05 83.858 ;
        RECT 79.76 77.082 91.769 77.139 ;
        RECT 85.004 71.838 85.05 83.858 ;
        RECT 73.008 83.834 85.004 83.904 ;
        RECT 79.806 77.036 91.815 77.093 ;
        RECT 84.958 71.884 85.004 83.904 ;
        RECT 72.962 83.88 84.958 83.95 ;
        RECT 79.852 76.99 91.861 77.047 ;
        RECT 84.912 71.93 84.958 83.95 ;
        RECT 72.916 83.926 84.912 83.996 ;
        RECT 79.898 76.944 110 77 ;
        RECT 84.866 71.976 84.912 83.996 ;
        RECT 72.87 83.972 84.866 84.042 ;
        RECT 79.944 76.898 110 77 ;
        RECT 84.82 72.022 84.866 84.042 ;
        RECT 72.824 84.018 84.82 84.088 ;
        RECT 79.99 76.852 110 77 ;
        RECT 84.774 72.068 84.82 84.088 ;
        RECT 72.778 84.064 84.774 84.134 ;
        RECT 80.036 76.806 110 77 ;
        RECT 84.728 72.114 84.774 84.134 ;
        RECT 72.732 84.11 84.728 84.18 ;
        RECT 80.082 76.76 110 77 ;
        RECT 84.682 72.16 84.728 84.18 ;
        RECT 72.686 84.156 84.682 84.226 ;
        RECT 80.128 76.714 110 77 ;
        RECT 84.636 72.206 84.682 84.226 ;
        RECT 72.64 84.202 84.636 84.272 ;
        RECT 80.174 76.668 110 77 ;
        RECT 84.59 72.252 84.636 84.272 ;
        RECT 72.594 84.248 84.59 84.318 ;
        RECT 80.22 76.622 110 77 ;
        RECT 84.544 72.298 84.59 84.318 ;
        RECT 72.548 84.294 84.544 84.364 ;
        RECT 80.266 76.576 110 77 ;
        RECT 84.498 72.344 84.544 84.364 ;
        RECT 72.502 84.34 84.498 84.41 ;
        RECT 80.312 76.53 110 77 ;
        RECT 84.452 72.39 84.498 84.41 ;
        RECT 72.456 84.386 84.452 84.456 ;
        RECT 80.358 76.484 110 77 ;
        RECT 84.406 72.436 84.452 84.456 ;
        RECT 72.41 84.432 84.406 84.502 ;
        RECT 80.404 76.438 110 77 ;
        RECT 84.36 72.482 84.406 84.502 ;
        RECT 72.364 84.478 84.36 84.548 ;
        RECT 80.45 76.392 110 77 ;
        RECT 84.314 72.528 84.36 84.548 ;
        RECT 72.318 84.524 84.314 84.594 ;
        RECT 80.496 76.346 110 77 ;
        RECT 84.268 72.574 84.314 84.594 ;
        RECT 72.272 84.57 84.268 84.64 ;
        RECT 80.542 76.3 110 77 ;
        RECT 84.222 72.62 84.268 84.64 ;
        RECT 72.226 84.616 84.222 84.686 ;
        RECT 80.588 76.254 110 77 ;
        RECT 84.176 72.666 84.222 84.686 ;
        RECT 72.18 84.662 84.176 84.732 ;
        RECT 80.634 76.208 110 77 ;
        RECT 84.13 72.712 84.176 84.732 ;
        RECT 72.134 84.708 84.13 84.778 ;
        RECT 80.68 76.162 110 77 ;
        RECT 84.084 72.758 84.13 84.778 ;
        RECT 72.088 84.754 84.084 84.824 ;
        RECT 80.726 76.116 110 77 ;
        RECT 84.038 72.804 84.084 84.824 ;
        RECT 72.042 84.8 84.038 84.87 ;
        RECT 80.772 76.07 110 77 ;
        RECT 83.992 72.85 84.038 84.87 ;
        RECT 71.996 84.846 83.992 84.916 ;
        RECT 80.818 76.024 110 77 ;
        RECT 83.946 72.896 83.992 84.916 ;
        RECT 71.95 84.892 83.946 84.962 ;
        RECT 80.864 75.978 110 77 ;
        RECT 83.9 72.942 83.946 84.962 ;
        RECT 71.904 84.938 83.9 85.008 ;
        RECT 80.91 75.932 110 77 ;
        RECT 83.854 72.988 83.9 85.008 ;
        RECT 71.858 84.984 83.854 85.054 ;
        RECT 80.956 75.886 110 77 ;
        RECT 83.808 73.034 83.854 85.054 ;
        RECT 71.812 85.03 83.808 85.1 ;
        RECT 81.002 75.84 110 77 ;
        RECT 83.762 73.08 83.808 85.1 ;
        RECT 71.766 85.076 83.762 85.146 ;
        RECT 81.048 75.794 110 77 ;
        RECT 83.716 73.126 83.762 85.146 ;
        RECT 71.72 85.122 83.716 85.192 ;
        RECT 81.094 75.748 110 77 ;
        RECT 83.67 73.172 83.716 85.192 ;
        RECT 71.674 85.168 83.67 85.238 ;
        RECT 81.14 75.702 110 77 ;
        RECT 83.624 73.218 83.67 85.238 ;
        RECT 71.628 85.214 83.624 85.284 ;
        RECT 81.186 75.656 110 77 ;
        RECT 83.578 73.264 83.624 85.284 ;
        RECT 71.582 85.26 83.578 85.33 ;
        RECT 81.232 75.61 110 77 ;
        RECT 83.532 73.31 83.578 85.33 ;
        RECT 71.536 85.306 83.532 85.376 ;
        RECT 81.278 75.564 110 77 ;
        RECT 83.486 73.356 83.532 85.376 ;
        RECT 71.49 85.352 83.486 85.422 ;
        RECT 81.324 75.518 110 77 ;
        RECT 83.44 73.402 83.486 85.422 ;
        RECT 71.444 85.398 83.44 85.468 ;
        RECT 81.37 75.472 110 77 ;
        RECT 83.394 73.448 83.44 85.468 ;
        RECT 71.398 85.444 83.394 85.514 ;
        RECT 81.416 75.426 110 77 ;
        RECT 83.348 73.494 83.394 85.514 ;
        RECT 71.352 85.49 83.348 85.56 ;
        RECT 81.462 75.38 110 77 ;
        RECT 83.302 73.54 83.348 85.56 ;
        RECT 71.306 85.536 83.302 85.606 ;
        RECT 81.508 75.334 110 77 ;
        RECT 83.256 73.586 83.302 85.606 ;
        RECT 71.26 85.582 83.256 85.652 ;
        RECT 81.554 75.288 110 77 ;
        RECT 83.21 73.632 83.256 85.652 ;
        RECT 71.214 85.628 83.21 85.698 ;
        RECT 81.6 75.242 110 77 ;
        RECT 83.164 73.678 83.21 85.698 ;
        RECT 71.168 85.674 83.164 85.744 ;
        RECT 81.646 75.196 110 77 ;
        RECT 83.118 73.724 83.164 85.744 ;
        RECT 71.122 85.72 83.118 85.79 ;
        RECT 81.692 75.15 110 77 ;
        RECT 83.072 73.77 83.118 85.79 ;
        RECT 71.076 85.766 83.072 85.836 ;
        RECT 81.738 75.104 110 77 ;
        RECT 83.026 73.816 83.072 85.836 ;
        RECT 71.03 85.812 83.026 85.882 ;
        RECT 81.784 75.058 110 77 ;
        RECT 82.98 73.862 83.026 85.882 ;
        RECT 70.984 85.858 82.98 85.928 ;
        RECT 81.83 75.012 110 77 ;
        RECT 82.934 73.908 82.98 85.928 ;
        RECT 70.938 85.904 82.934 85.974 ;
        RECT 81.876 74.966 110 77 ;
        RECT 82.888 73.954 82.934 85.974 ;
        RECT 70.892 85.95 82.888 86.02 ;
        RECT 81.922 74.92 110 77 ;
        RECT 82.842 74 82.888 86.02 ;
        RECT 70.846 85.996 82.842 86.066 ;
        RECT 81.968 74.874 110 77 ;
        RECT 82.796 74.046 82.842 86.066 ;
        RECT 70.8 86.042 82.796 86.112 ;
        RECT 82.014 74.828 110 77 ;
        RECT 82.75 74.092 82.796 86.112 ;
        RECT 70.754 86.088 82.75 86.158 ;
        RECT 82.06 74.782 110 77 ;
        RECT 82.704 74.138 82.75 86.158 ;
        RECT 70.708 86.134 82.704 86.204 ;
        RECT 82.106 74.736 110 77 ;
        RECT 82.658 74.184 82.704 86.204 ;
        RECT 70.662 86.18 82.658 86.25 ;
        RECT 82.152 74.69 110 77 ;
        RECT 82.612 74.23 82.658 86.25 ;
        RECT 70.616 86.226 82.612 86.296 ;
        RECT 82.198 74.644 110 77 ;
        RECT 82.566 74.276 82.612 86.296 ;
        RECT 70.57 86.272 82.566 86.342 ;
        RECT 82.244 74.598 110 77 ;
        RECT 82.52 74.322 82.566 86.342 ;
        RECT 70.524 86.318 82.52 86.388 ;
        RECT 82.29 74.552 110 77 ;
        RECT 82.474 74.368 82.52 86.388 ;
        RECT 70.478 86.364 82.474 86.434 ;
        RECT 82.336 74.506 110 77 ;
        RECT 82.428 74.414 82.474 86.434 ;
        RECT 70.432 86.41 82.428 86.48 ;
        RECT 82.382 74.46 110 77 ;
        RECT 70.386 86.456 82.382 86.526 ;
        RECT 70.34 86.502 82.336 86.572 ;
        RECT 70.294 86.548 82.29 86.618 ;
        RECT 70.248 86.594 82.244 86.664 ;
        RECT 70.202 86.64 82.198 86.71 ;
        RECT 70.156 86.686 82.152 86.756 ;
        RECT 70.11 86.732 82.106 86.802 ;
        RECT 70.064 86.778 82.06 86.848 ;
        RECT 70.018 86.824 82.014 86.894 ;
        RECT 69.972 86.87 81.968 86.94 ;
        RECT 69.926 86.916 81.922 86.986 ;
        RECT 69.88 86.962 81.876 87.032 ;
        RECT 69.834 87.008 81.83 87.078 ;
        RECT 69.788 87.054 81.784 87.124 ;
        RECT 69.742 87.1 81.738 87.17 ;
        RECT 69.696 87.146 81.692 87.216 ;
        RECT 69.65 87.192 81.646 87.262 ;
        RECT 69.604 87.238 81.6 87.308 ;
        RECT 69.558 87.284 81.554 87.354 ;
        RECT 69.512 87.33 81.508 87.4 ;
        RECT 69.466 87.376 81.462 87.446 ;
        RECT 69.42 87.422 81.416 87.492 ;
        RECT 69.374 87.468 81.37 87.538 ;
        RECT 69.328 87.514 81.324 87.584 ;
        RECT 69.282 87.56 81.278 87.63 ;
        RECT 69.236 87.606 81.232 87.676 ;
        RECT 69.19 87.652 81.186 87.722 ;
        RECT 69.144 87.698 81.14 87.768 ;
        RECT 69.098 87.744 81.094 87.814 ;
        RECT 69.052 87.79 81.048 87.86 ;
        RECT 69.006 87.836 81.002 87.906 ;
        RECT 68.96 87.882 80.956 87.952 ;
        RECT 68.914 87.928 80.91 87.998 ;
        RECT 68.868 87.974 80.864 88.044 ;
        RECT 68.822 88.02 80.818 88.09 ;
        RECT 68.776 88.066 80.772 88.136 ;
        RECT 68.73 88.112 80.726 88.182 ;
        RECT 68.684 88.158 80.68 88.228 ;
        RECT 68.638 88.204 80.634 88.274 ;
        RECT 68.592 88.25 80.588 88.32 ;
        RECT 68.546 88.296 80.542 88.366 ;
        RECT 68.5 88.342 80.496 88.412 ;
        RECT 68.5 88.342 80.45 88.458 ;
        RECT 68.5 88.342 80.404 88.504 ;
        RECT 68.5 88.342 80.358 88.55 ;
        RECT 68.5 88.342 80.312 88.596 ;
        RECT 68.5 88.342 80.266 88.642 ;
        RECT 68.5 88.342 80.22 88.688 ;
        RECT 68.5 88.342 80.174 88.734 ;
        RECT 68.5 88.342 80.128 88.78 ;
        RECT 68.5 88.342 80.082 88.826 ;
        RECT 68.5 88.342 80.036 88.872 ;
        RECT 68.5 88.342 79.99 88.918 ;
        RECT 68.5 88.342 79.944 88.964 ;
        RECT 68.5 88.342 79.898 89.01 ;
        RECT 68.5 88.342 79.852 89.056 ;
        RECT 68.5 88.342 79.806 89.102 ;
        RECT 68.5 88.342 79.76 89.148 ;
        RECT 68.5 88.342 79.714 89.194 ;
        RECT 68.5 88.342 79.668 89.24 ;
        RECT 68.5 88.342 79.622 89.286 ;
        RECT 68.5 88.342 79.576 89.332 ;
        RECT 68.5 88.342 79.53 89.378 ;
        RECT 68.5 88.342 79.484 89.424 ;
        RECT 68.5 88.342 79.438 89.47 ;
        RECT 68.5 88.342 79.392 89.516 ;
        RECT 68.5 88.342 79.346 89.562 ;
        RECT 68.5 88.342 79.3 89.608 ;
        RECT 68.5 88.342 79.254 89.654 ;
        RECT 68.5 88.342 79.208 89.7 ;
        RECT 68.5 88.342 79.162 89.746 ;
        RECT 68.5 88.342 79.116 89.792 ;
        RECT 68.5 88.342 79.07 89.838 ;
        RECT 68.5 88.342 79.024 89.884 ;
        RECT 68.5 88.342 78.978 89.93 ;
        RECT 68.5 88.342 78.932 89.976 ;
        RECT 68.5 88.342 78.886 90.022 ;
        RECT 68.5 88.342 78.84 90.068 ;
        RECT 68.5 88.342 78.794 90.114 ;
        RECT 68.5 88.342 78.748 90.16 ;
        RECT 68.5 88.342 78.702 90.206 ;
        RECT 68.5 88.342 78.656 90.252 ;
        RECT 68.5 88.342 78.61 90.298 ;
        RECT 68.5 88.342 78.564 90.344 ;
        RECT 68.5 88.342 78.518 90.39 ;
        RECT 68.5 88.342 78.472 90.436 ;
        RECT 68.5 88.342 78.426 90.482 ;
        RECT 68.5 88.342 78.38 90.528 ;
        RECT 68.5 88.342 78.334 90.574 ;
        RECT 68.5 88.342 78.288 90.62 ;
        RECT 68.5 88.342 78.242 90.666 ;
        RECT 68.5 88.342 78.196 90.712 ;
        RECT 68.5 88.342 78.15 90.758 ;
        RECT 68.5 88.342 78.104 90.804 ;
        RECT 68.5 88.342 78.058 90.85 ;
        RECT 68.5 88.342 78.012 90.896 ;
        RECT 68.5 88.342 77.966 90.942 ;
        RECT 68.5 88.342 77.92 90.988 ;
        RECT 68.5 88.342 77.874 91.034 ;
        RECT 68.5 88.342 77.828 91.08 ;
        RECT 68.5 88.342 77.782 91.126 ;
        RECT 68.5 88.342 77.736 91.172 ;
        RECT 68.5 88.342 77.69 91.218 ;
        RECT 68.5 88.342 77.644 91.264 ;
        RECT 68.5 88.342 77.598 91.31 ;
        RECT 68.5 88.342 77.552 91.356 ;
        RECT 68.5 88.342 77.506 91.402 ;
        RECT 68.5 88.342 77.46 91.448 ;
        RECT 68.5 88.342 77.414 91.494 ;
        RECT 68.5 88.342 77.368 91.54 ;
        RECT 68.5 88.342 77.322 91.586 ;
        RECT 68.5 88.342 77.276 91.632 ;
        RECT 68.5 88.342 77.23 91.678 ;
        RECT 68.5 88.342 77.184 91.724 ;
        RECT 68.5 88.342 77.138 91.77 ;
        RECT 68.5 88.342 77.092 91.816 ;
        RECT 68.5 88.342 77.046 91.862 ;
        RECT 68.5 88.342 77 110 ;
        RECT 75.642 44.6 75.688 61.57 ;
        RECT 58.714 61.528 75.642 61.616 ;
        RECT 60.002 60.24 76.955 60.303 ;
        RECT 75.596 44.646 75.642 61.616 ;
        RECT 58.668 61.574 75.596 61.662 ;
        RECT 60.048 60.194 77.001 60.257 ;
        RECT 75.55 44.692 75.596 61.662 ;
        RECT 58.622 61.62 75.55 61.708 ;
        RECT 60.094 60.148 77.047 60.211 ;
        RECT 75.504 44.738 75.55 61.708 ;
        RECT 58.576 61.666 75.504 61.754 ;
        RECT 60.14 60.102 77.093 60.165 ;
        RECT 75.458 44.784 75.504 61.754 ;
        RECT 58.53 61.712 75.458 61.8 ;
        RECT 60.186 60.056 77.139 60.119 ;
        RECT 75.412 44.83 75.458 61.8 ;
        RECT 58.484 61.758 75.412 61.846 ;
        RECT 60.232 60.01 77.185 60.073 ;
        RECT 75.366 44.876 75.412 61.846 ;
        RECT 58.438 61.804 75.366 61.892 ;
        RECT 60.278 59.964 77.231 60.027 ;
        RECT 75.32 44.922 75.366 61.892 ;
        RECT 58.392 61.85 75.32 61.938 ;
        RECT 60.324 59.918 77.277 59.981 ;
        RECT 75.274 44.968 75.32 61.938 ;
        RECT 58.346 61.896 75.274 61.984 ;
        RECT 60.37 59.872 77.323 59.935 ;
        RECT 75.228 45.014 75.274 61.984 ;
        RECT 58.3 61.942 75.228 62.03 ;
        RECT 60.416 59.826 77.369 59.889 ;
        RECT 75.182 45.06 75.228 62.03 ;
        RECT 58.254 61.988 75.182 62.076 ;
        RECT 60.462 59.78 77.415 59.843 ;
        RECT 75.136 45.106 75.182 62.076 ;
        RECT 58.208 62.034 75.136 62.122 ;
        RECT 60.508 59.734 77.461 59.797 ;
        RECT 75.09 45.152 75.136 62.122 ;
        RECT 58.162 62.08 75.09 62.168 ;
        RECT 60.554 59.688 77.507 59.751 ;
        RECT 75.044 45.198 75.09 62.168 ;
        RECT 58.116 62.126 75.044 62.214 ;
        RECT 60.6 59.642 77.553 59.705 ;
        RECT 74.998 45.244 75.044 62.214 ;
        RECT 58.07 62.172 74.998 62.26 ;
        RECT 60.646 59.596 77.599 59.659 ;
        RECT 74.952 45.29 74.998 62.26 ;
        RECT 58.024 62.218 74.952 62.306 ;
        RECT 60.692 59.55 77.645 59.613 ;
        RECT 74.906 45.336 74.952 62.306 ;
        RECT 57.978 62.264 74.906 62.352 ;
        RECT 60.738 59.504 77.691 59.567 ;
        RECT 74.86 45.382 74.906 62.352 ;
        RECT 57.932 62.31 74.86 62.398 ;
        RECT 60.784 59.458 77.737 59.521 ;
        RECT 74.814 45.428 74.86 62.398 ;
        RECT 57.886 62.356 74.814 62.444 ;
        RECT 60.83 59.412 77.783 59.475 ;
        RECT 74.768 45.474 74.814 62.444 ;
        RECT 57.84 62.402 74.768 62.49 ;
        RECT 60.876 59.366 77.829 59.429 ;
        RECT 74.722 45.52 74.768 62.49 ;
        RECT 57.794 62.448 74.722 62.536 ;
        RECT 60.922 59.32 77.875 59.383 ;
        RECT 74.676 45.566 74.722 62.536 ;
        RECT 57.748 62.494 74.676 62.582 ;
        RECT 60.968 59.274 77.921 59.337 ;
        RECT 74.63 45.612 74.676 62.582 ;
        RECT 57.702 62.54 74.63 62.628 ;
        RECT 61.014 59.228 77.967 59.291 ;
        RECT 74.584 45.658 74.63 62.628 ;
        RECT 57.656 62.586 74.584 62.674 ;
        RECT 61.06 59.182 78.013 59.245 ;
        RECT 74.538 45.704 74.584 62.674 ;
        RECT 57.61 62.632 74.538 62.72 ;
        RECT 61.106 59.136 78.059 59.199 ;
        RECT 74.492 45.75 74.538 62.72 ;
        RECT 57.564 62.678 74.492 62.766 ;
        RECT 61.152 59.09 78.105 59.153 ;
        RECT 74.446 45.796 74.492 62.766 ;
        RECT 57.518 62.724 74.446 62.812 ;
        RECT 61.198 59.044 78.151 59.107 ;
        RECT 74.4 45.842 74.446 62.812 ;
        RECT 57.472 62.77 74.4 62.858 ;
        RECT 61.244 58.998 78.197 59.061 ;
        RECT 74.354 45.888 74.4 62.858 ;
        RECT 57.426 62.816 74.354 62.904 ;
        RECT 61.29 58.952 78.243 59.015 ;
        RECT 74.308 45.934 74.354 62.904 ;
        RECT 57.38 62.862 74.308 62.95 ;
        RECT 61.336 58.906 78.289 58.969 ;
        RECT 74.262 45.98 74.308 62.95 ;
        RECT 57.334 62.908 74.262 62.996 ;
        RECT 61.382 58.86 78.335 58.923 ;
        RECT 74.216 46.026 74.262 62.996 ;
        RECT 57.288 62.954 74.216 63.042 ;
        RECT 61.428 58.814 78.381 58.877 ;
        RECT 74.17 46.072 74.216 63.042 ;
        RECT 57.242 63 74.17 63.088 ;
        RECT 61.474 58.768 78.427 58.831 ;
        RECT 74.124 46.118 74.17 63.088 ;
        RECT 57.196 63.046 74.124 63.134 ;
        RECT 61.52 58.722 78.473 58.785 ;
        RECT 74.078 46.164 74.124 63.134 ;
        RECT 57.15 63.092 74.078 63.18 ;
        RECT 61.566 58.676 78.519 58.739 ;
        RECT 74.032 46.21 74.078 63.18 ;
        RECT 57.104 63.138 74.032 63.226 ;
        RECT 61.612 58.63 78.565 58.693 ;
        RECT 73.986 46.256 74.032 63.226 ;
        RECT 57.058 63.184 73.986 63.272 ;
        RECT 61.658 58.584 78.611 58.647 ;
        RECT 73.94 46.302 73.986 63.272 ;
        RECT 57.012 63.23 73.94 63.318 ;
        RECT 61.704 58.538 78.657 58.601 ;
        RECT 73.894 46.348 73.94 63.318 ;
        RECT 56.966 63.276 73.894 63.364 ;
        RECT 61.75 58.492 78.703 58.555 ;
        RECT 73.848 46.394 73.894 63.364 ;
        RECT 56.92 63.322 73.848 63.41 ;
        RECT 61.796 58.446 78.749 58.509 ;
        RECT 73.802 46.44 73.848 63.41 ;
        RECT 56.874 63.368 73.802 63.456 ;
        RECT 61.842 58.4 78.795 58.463 ;
        RECT 73.756 46.486 73.802 63.456 ;
        RECT 56.828 63.414 73.756 63.502 ;
        RECT 61.888 58.354 78.841 58.417 ;
        RECT 73.71 46.532 73.756 63.502 ;
        RECT 56.782 63.46 73.71 63.548 ;
        RECT 61.934 58.308 78.887 58.371 ;
        RECT 73.664 46.578 73.71 63.548 ;
        RECT 56.736 63.506 73.664 63.594 ;
        RECT 61.98 58.262 78.933 58.325 ;
        RECT 73.618 46.624 73.664 63.594 ;
        RECT 56.69 63.552 73.618 63.64 ;
        RECT 62.026 58.216 78.979 58.279 ;
        RECT 73.572 46.67 73.618 63.64 ;
        RECT 56.644 63.598 73.572 63.686 ;
        RECT 62.072 58.17 79.025 58.233 ;
        RECT 73.526 46.716 73.572 63.686 ;
        RECT 56.598 63.644 73.526 63.732 ;
        RECT 62.118 58.124 79.071 58.187 ;
        RECT 73.48 46.762 73.526 63.732 ;
        RECT 56.552 63.69 73.48 63.778 ;
        RECT 62.164 58.078 79.117 58.141 ;
        RECT 73.434 46.808 73.48 63.778 ;
        RECT 56.506 63.736 73.434 63.824 ;
        RECT 62.21 58.032 79.163 58.095 ;
        RECT 73.388 46.854 73.434 63.824 ;
        RECT 56.46 63.782 73.388 63.87 ;
        RECT 62.256 57.986 79.209 58.049 ;
        RECT 73.342 46.9 73.388 63.87 ;
        RECT 56.414 63.828 73.342 63.916 ;
        RECT 62.302 57.94 79.255 58.003 ;
        RECT 73.296 46.946 73.342 63.916 ;
        RECT 56.368 63.874 73.296 63.962 ;
        RECT 62.348 57.894 79.301 57.957 ;
        RECT 73.25 46.992 73.296 63.962 ;
        RECT 56.322 63.92 73.25 64.008 ;
        RECT 62.394 57.848 79.347 57.911 ;
        RECT 73.204 47.038 73.25 64.008 ;
        RECT 56.276 63.966 73.204 64.054 ;
        RECT 62.44 57.802 79.393 57.865 ;
        RECT 73.158 47.084 73.204 64.054 ;
        RECT 56.23 64.012 73.158 64.1 ;
        RECT 62.486 57.756 79.439 57.819 ;
        RECT 73.112 47.13 73.158 64.1 ;
        RECT 56.184 64.058 73.112 64.146 ;
        RECT 62.532 57.71 79.485 57.773 ;
        RECT 73.066 47.176 73.112 64.146 ;
        RECT 56.138 64.104 73.066 64.192 ;
        RECT 62.578 57.664 79.531 57.727 ;
        RECT 73.02 47.222 73.066 64.192 ;
        RECT 56.092 64.15 73.02 64.238 ;
        RECT 62.624 57.618 79.577 57.681 ;
        RECT 72.974 47.268 73.02 64.238 ;
        RECT 56 64.242 72.974 64.284 ;
        RECT 56.046 64.196 72.974 64.284 ;
        RECT 62.67 57.572 79.623 57.635 ;
        RECT 72.928 47.314 72.974 64.284 ;
        RECT 55.96 64.285 72.928 64.33 ;
        RECT 62.716 57.526 79.669 57.589 ;
        RECT 72.882 47.36 72.928 64.33 ;
        RECT 55.914 64.328 72.882 64.376 ;
        RECT 62.762 57.48 79.715 57.543 ;
        RECT 72.836 47.406 72.882 64.376 ;
        RECT 55.868 64.374 72.836 64.422 ;
        RECT 62.808 57.434 79.761 57.497 ;
        RECT 72.79 47.452 72.836 64.422 ;
        RECT 55.822 64.42 72.79 64.468 ;
        RECT 62.854 57.388 79.807 57.451 ;
        RECT 72.744 47.498 72.79 64.468 ;
        RECT 55.776 64.466 72.744 64.514 ;
        RECT 62.9 57.342 79.853 57.405 ;
        RECT 72.698 47.544 72.744 64.514 ;
        RECT 55.73 64.512 72.698 64.56 ;
        RECT 62.946 57.296 79.899 57.359 ;
        RECT 72.652 47.59 72.698 64.56 ;
        RECT 55.684 64.558 72.652 64.606 ;
        RECT 62.992 57.25 79.945 57.313 ;
        RECT 72.606 47.636 72.652 64.606 ;
        RECT 55.638 64.604 72.606 64.652 ;
        RECT 63.038 57.204 79.991 57.267 ;
        RECT 72.56 47.682 72.606 64.652 ;
        RECT 55.592 64.65 72.56 64.698 ;
        RECT 63.084 57.158 80.037 57.221 ;
        RECT 72.514 47.728 72.56 64.698 ;
        RECT 55.546 64.696 72.514 64.744 ;
        RECT 63.13 57.112 80.083 57.175 ;
        RECT 72.468 47.774 72.514 64.744 ;
        RECT 55.5 64.742 72.468 64.79 ;
        RECT 63.176 57.066 80.129 57.129 ;
        RECT 72.422 47.82 72.468 64.79 ;
        RECT 55.454 64.788 72.422 64.836 ;
        RECT 63.222 57.02 80.175 57.083 ;
        RECT 72.376 47.866 72.422 64.836 ;
        RECT 55.408 64.834 72.376 64.882 ;
        RECT 63.268 56.974 80.221 57.037 ;
        RECT 72.33 47.912 72.376 64.882 ;
        RECT 55.362 64.88 72.33 64.928 ;
        RECT 63.314 56.928 80.267 56.991 ;
        RECT 72.284 47.958 72.33 64.928 ;
        RECT 55.316 64.926 72.284 64.974 ;
        RECT 63.36 56.882 80.313 56.945 ;
        RECT 72.238 48.004 72.284 64.974 ;
        RECT 55.27 64.972 72.238 65.02 ;
        RECT 63.406 56.836 80.359 56.899 ;
        RECT 72.192 48.05 72.238 65.02 ;
        RECT 55.224 65.018 72.192 65.066 ;
        RECT 63.452 56.79 80.405 56.853 ;
        RECT 72.146 48.096 72.192 65.066 ;
        RECT 55.178 65.064 72.146 65.112 ;
        RECT 63.498 56.744 80.451 56.807 ;
        RECT 72.1 48.142 72.146 65.112 ;
        RECT 55.132 65.11 72.1 65.158 ;
        RECT 63.544 56.698 80.497 56.761 ;
        RECT 72.054 48.188 72.1 65.158 ;
        RECT 55.086 65.156 72.054 65.204 ;
        RECT 63.59 56.652 80.543 56.715 ;
        RECT 72.008 48.234 72.054 65.204 ;
        RECT 55.04 65.202 72.008 65.25 ;
        RECT 63.636 56.606 80.589 56.669 ;
        RECT 71.962 48.28 72.008 65.25 ;
        RECT 54.994 65.248 71.962 65.296 ;
        RECT 63.682 56.56 80.635 56.623 ;
        RECT 71.916 48.326 71.962 65.296 ;
        RECT 54.948 65.294 71.916 65.342 ;
        RECT 63.728 56.514 80.681 56.577 ;
        RECT 71.87 48.372 71.916 65.342 ;
        RECT 54.902 65.34 71.87 65.388 ;
        RECT 63.774 56.468 80.727 56.531 ;
        RECT 71.824 48.418 71.87 65.388 ;
        RECT 54.856 65.386 71.824 65.434 ;
        RECT 63.82 56.422 80.773 56.485 ;
        RECT 71.778 48.464 71.824 65.434 ;
        RECT 54.81 65.432 71.778 65.48 ;
        RECT 63.866 56.376 80.819 56.439 ;
        RECT 71.732 48.51 71.778 65.48 ;
        RECT 54.764 65.478 71.732 65.526 ;
        RECT 63.912 56.33 80.865 56.393 ;
        RECT 71.686 48.556 71.732 65.526 ;
        RECT 54.718 65.524 71.686 65.572 ;
        RECT 63.958 56.284 80.911 56.347 ;
        RECT 71.64 48.602 71.686 65.572 ;
        RECT 54.672 65.57 71.64 65.618 ;
        RECT 64.004 56.238 80.957 56.301 ;
        RECT 71.594 48.648 71.64 65.618 ;
        RECT 54.626 65.616 71.594 65.664 ;
        RECT 64.05 56.192 81.003 56.255 ;
        RECT 71.548 48.694 71.594 65.664 ;
        RECT 54.58 65.662 71.548 65.71 ;
        RECT 64.096 56.146 81.049 56.209 ;
        RECT 71.502 48.74 71.548 65.71 ;
        RECT 54.534 65.708 71.502 65.756 ;
        RECT 64.142 56.1 81.095 56.163 ;
        RECT 71.456 48.786 71.502 65.756 ;
        RECT 54.488 65.754 71.456 65.802 ;
        RECT 64.188 56.054 81.141 56.117 ;
        RECT 71.41 48.832 71.456 65.802 ;
        RECT 54.442 65.8 71.41 65.848 ;
        RECT 64.234 56.008 81.187 56.071 ;
        RECT 71.364 48.878 71.41 65.848 ;
        RECT 54.396 65.846 71.364 65.894 ;
        RECT 64.28 55.962 81.233 56.024 ;
        RECT 71.318 48.924 71.364 65.894 ;
        RECT 54.35 65.892 71.318 65.94 ;
        RECT 64.326 55.916 110 56 ;
        RECT 71.272 48.97 71.318 65.94 ;
        RECT 54.304 65.938 71.272 65.986 ;
        RECT 64.372 55.87 110 56 ;
        RECT 71.226 49.016 71.272 65.986 ;
        RECT 54.258 65.984 71.226 66.032 ;
        RECT 64.418 55.824 110 56 ;
        RECT 71.18 49.062 71.226 66.032 ;
        RECT 54.212 66.03 71.18 66.078 ;
        RECT 64.464 55.778 110 56 ;
        RECT 71.134 49.108 71.18 66.078 ;
        RECT 54.166 66.076 71.134 66.124 ;
        RECT 64.51 55.732 110 56 ;
        RECT 71.088 49.154 71.134 66.124 ;
        RECT 54.12 66.122 71.088 66.17 ;
        RECT 64.556 55.686 110 56 ;
        RECT 71.042 49.2 71.088 66.17 ;
        RECT 54.074 66.168 71.042 66.216 ;
        RECT 64.602 55.64 110 56 ;
        RECT 70.996 49.246 71.042 66.216 ;
        RECT 54.028 66.214 70.996 66.262 ;
        RECT 64.648 55.594 110 56 ;
        RECT 70.95 49.292 70.996 66.262 ;
        RECT 53.982 66.26 70.95 66.308 ;
        RECT 64.694 55.548 110 56 ;
        RECT 70.904 49.338 70.95 66.308 ;
        RECT 53.936 66.306 70.904 66.354 ;
        RECT 64.74 55.502 110 56 ;
        RECT 70.858 49.384 70.904 66.354 ;
        RECT 53.89 66.352 70.858 66.4 ;
        RECT 64.786 55.456 110 56 ;
        RECT 70.812 49.43 70.858 66.4 ;
        RECT 53.844 66.398 70.812 66.446 ;
        RECT 64.832 55.41 110 56 ;
        RECT 70.766 49.476 70.812 66.446 ;
        RECT 53.798 66.444 70.766 66.492 ;
        RECT 64.878 55.364 110 56 ;
        RECT 70.72 49.522 70.766 66.492 ;
        RECT 53.752 66.49 70.72 66.538 ;
        RECT 64.924 55.318 110 56 ;
        RECT 70.674 49.568 70.72 66.538 ;
        RECT 53.706 66.536 70.674 66.584 ;
        RECT 64.97 55.272 110 56 ;
        RECT 70.628 49.614 70.674 66.584 ;
        RECT 53.66 66.582 70.628 66.63 ;
        RECT 65.016 55.226 110 56 ;
        RECT 70.582 49.66 70.628 66.63 ;
        RECT 53.614 66.628 70.582 66.676 ;
        RECT 65.062 55.18 110 56 ;
        RECT 70.536 49.706 70.582 66.676 ;
        RECT 53.568 66.674 70.536 66.722 ;
        RECT 65.108 55.134 110 56 ;
        RECT 70.49 49.752 70.536 66.722 ;
        RECT 53.522 66.72 70.49 66.768 ;
        RECT 65.154 55.088 110 56 ;
        RECT 70.444 49.798 70.49 66.768 ;
        RECT 53.476 66.766 70.444 66.814 ;
        RECT 65.2 55.042 110 56 ;
        RECT 70.398 49.844 70.444 66.814 ;
        RECT 53.43 66.812 70.398 66.86 ;
        RECT 65.246 54.996 110 56 ;
        RECT 70.352 49.89 70.398 66.86 ;
        RECT 53.384 66.858 70.352 66.906 ;
        RECT 65.292 54.95 110 56 ;
        RECT 70.306 49.936 70.352 66.906 ;
        RECT 53.338 66.904 70.306 66.952 ;
        RECT 65.338 54.904 110 56 ;
        RECT 70.26 49.982 70.306 66.952 ;
        RECT 53.292 66.95 70.26 66.998 ;
        RECT 65.384 54.858 110 56 ;
        RECT 70.214 50.028 70.26 66.998 ;
        RECT 53.246 66.996 70.214 67.044 ;
        RECT 65.43 54.812 110 56 ;
        RECT 70.168 50.074 70.214 67.044 ;
        RECT 53.2 67.042 70.168 67.09 ;
        RECT 65.476 54.766 110 56 ;
        RECT 70.122 50.12 70.168 67.09 ;
        RECT 53.154 67.088 70.122 67.136 ;
        RECT 65.522 54.72 110 56 ;
        RECT 70.076 50.166 70.122 67.136 ;
        RECT 53.108 67.134 70.076 67.182 ;
        RECT 65.568 54.674 110 56 ;
        RECT 70.03 50.212 70.076 67.182 ;
        RECT 53.062 67.18 70.03 67.228 ;
        RECT 65.614 54.628 110 56 ;
        RECT 69.984 50.258 70.03 67.228 ;
        RECT 53.016 67.226 69.984 67.274 ;
        RECT 65.66 54.582 110 56 ;
        RECT 69.938 50.304 69.984 67.274 ;
        RECT 52.97 67.272 69.938 67.32 ;
        RECT 65.706 54.536 110 56 ;
        RECT 69.892 50.35 69.938 67.32 ;
        RECT 52.924 67.318 69.892 67.366 ;
        RECT 65.752 54.49 110 56 ;
        RECT 69.846 50.396 69.892 67.366 ;
        RECT 52.878 67.364 69.846 67.412 ;
        RECT 65.798 54.444 110 56 ;
        RECT 69.8 50.442 69.846 67.412 ;
        RECT 52.832 67.41 69.8 67.458 ;
        RECT 65.844 54.398 110 56 ;
        RECT 69.754 50.488 69.8 67.458 ;
        RECT 52.786 67.456 69.754 67.504 ;
        RECT 65.89 54.352 110 56 ;
        RECT 69.708 50.534 69.754 67.504 ;
        RECT 52.74 67.502 69.708 67.55 ;
        RECT 65.936 54.306 110 56 ;
        RECT 69.662 50.58 69.708 67.55 ;
        RECT 52.694 67.548 69.662 67.596 ;
        RECT 65.982 54.26 110 56 ;
        RECT 69.616 50.626 69.662 67.596 ;
        RECT 52.648 67.594 69.616 67.642 ;
        RECT 66.028 54.214 110 56 ;
        RECT 69.57 50.672 69.616 67.642 ;
        RECT 52.602 67.64 69.57 67.688 ;
        RECT 66.074 54.168 110 56 ;
        RECT 69.524 50.718 69.57 67.688 ;
        RECT 52.556 67.686 69.524 67.734 ;
        RECT 66.12 54.122 110 56 ;
        RECT 69.478 50.764 69.524 67.734 ;
        RECT 52.51 67.732 69.478 67.78 ;
        RECT 66.166 54.076 110 56 ;
        RECT 69.432 50.81 69.478 67.78 ;
        RECT 52.464 67.778 69.432 67.826 ;
        RECT 66.212 54.03 110 56 ;
        RECT 69.386 50.856 69.432 67.826 ;
        RECT 52.418 67.824 69.386 67.872 ;
        RECT 66.258 53.984 110 56 ;
        RECT 69.34 50.902 69.386 67.872 ;
        RECT 52.372 67.87 69.34 67.918 ;
        RECT 66.304 53.938 110 56 ;
        RECT 69.294 50.948 69.34 67.918 ;
        RECT 52.326 67.916 69.294 67.964 ;
        RECT 66.35 53.892 110 56 ;
        RECT 69.248 50.994 69.294 67.964 ;
        RECT 52.28 67.962 69.248 68.01 ;
        RECT 66.396 53.846 110 56 ;
        RECT 69.202 51.04 69.248 68.01 ;
        RECT 52.234 68.008 69.202 68.056 ;
        RECT 66.442 53.8 110 56 ;
        RECT 69.156 51.086 69.202 68.056 ;
        RECT 52.188 68.054 69.156 68.102 ;
        RECT 66.488 53.754 110 56 ;
        RECT 69.11 51.132 69.156 68.102 ;
        RECT 52.142 68.1 69.11 68.148 ;
        RECT 66.534 53.708 110 56 ;
        RECT 69.064 51.178 69.11 68.148 ;
        RECT 52.096 68.146 69.064 68.194 ;
        RECT 66.58 53.662 110 56 ;
        RECT 69.018 51.224 69.064 68.194 ;
        RECT 52.05 68.192 69.018 68.24 ;
        RECT 66.626 53.616 110 56 ;
        RECT 68.972 51.27 69.018 68.24 ;
        RECT 52.004 68.238 68.972 68.286 ;
        RECT 66.672 53.57 110 56 ;
        RECT 68.926 51.316 68.972 68.286 ;
        RECT 51.958 68.284 68.926 68.332 ;
        RECT 66.718 53.524 110 56 ;
        RECT 68.88 51.362 68.926 68.332 ;
        RECT 51.912 68.33 68.88 68.378 ;
        RECT 66.764 53.478 110 56 ;
        RECT 68.834 51.408 68.88 68.378 ;
        RECT 51.866 68.376 68.834 68.424 ;
        RECT 66.81 53.432 110 56 ;
        RECT 68.788 51.454 68.834 68.424 ;
        RECT 51.82 68.422 68.788 68.47 ;
        RECT 66.856 53.386 110 56 ;
        RECT 68.742 51.5 68.788 68.47 ;
        RECT 51.774 68.468 68.742 68.516 ;
        RECT 66.902 53.34 110 56 ;
        RECT 68.696 51.546 68.742 68.516 ;
        RECT 51.728 68.514 68.696 68.562 ;
        RECT 66.948 53.294 110 56 ;
        RECT 68.65 51.592 68.696 68.562 ;
        RECT 51.682 68.56 68.65 68.608 ;
        RECT 66.994 53.248 110 56 ;
        RECT 68.604 51.638 68.65 68.608 ;
        RECT 51.636 68.606 68.604 68.654 ;
        RECT 67.04 53.202 110 56 ;
        RECT 68.558 51.684 68.604 68.654 ;
        RECT 51.59 68.652 68.558 68.7 ;
        RECT 67.086 53.156 110 56 ;
        RECT 68.512 51.73 68.558 68.7 ;
        RECT 51.544 68.698 68.512 68.746 ;
        RECT 67.132 53.11 110 56 ;
        RECT 68.466 51.776 68.512 68.746 ;
        RECT 51.498 68.744 68.466 68.792 ;
        RECT 67.178 53.064 110 56 ;
        RECT 68.42 51.822 68.466 68.792 ;
        RECT 51.452 68.79 68.42 68.838 ;
        RECT 67.224 53.018 110 56 ;
        RECT 68.374 51.868 68.42 68.838 ;
        RECT 51.406 68.836 68.374 68.884 ;
        RECT 67.27 52.972 110 56 ;
        RECT 68.328 51.914 68.374 68.884 ;
        RECT 51.36 68.882 68.328 68.93 ;
        RECT 67.316 52.926 110 56 ;
        RECT 68.282 51.96 68.328 68.93 ;
        RECT 51.314 68.928 68.282 68.976 ;
        RECT 67.362 52.88 110 56 ;
        RECT 68.236 52.006 68.282 68.976 ;
        RECT 51.268 68.974 68.236 69.022 ;
        RECT 67.408 52.834 110 56 ;
        RECT 68.19 52.052 68.236 69.022 ;
        RECT 51.222 69.02 68.19 69.068 ;
        RECT 67.454 52.788 110 56 ;
        RECT 68.144 52.098 68.19 69.068 ;
        RECT 51.176 69.066 68.144 69.114 ;
        RECT 67.5 52.742 110 56 ;
        RECT 68.098 52.144 68.144 69.114 ;
        RECT 51.13 69.112 68.098 69.16 ;
        RECT 67.546 52.696 110 56 ;
        RECT 68.052 52.19 68.098 69.16 ;
        RECT 51.084 69.158 68.052 69.206 ;
        RECT 67.592 52.65 110 56 ;
        RECT 68.006 52.236 68.052 69.206 ;
        RECT 51.038 69.204 68.006 69.252 ;
        RECT 67.638 52.604 110 56 ;
        RECT 67.96 52.282 68.006 69.252 ;
        RECT 50.992 69.25 67.96 69.298 ;
        RECT 67.684 52.558 110 56 ;
        RECT 67.914 52.328 67.96 69.298 ;
        RECT 50.946 69.296 67.914 69.344 ;
        RECT 67.73 52.512 110 56 ;
        RECT 67.868 52.374 67.914 69.344 ;
        RECT 50.9 69.342 67.868 69.39 ;
        RECT 67.776 52.466 110 56 ;
        RECT 67.822 52.42 67.868 69.39 ;
        RECT 50.854 69.388 67.822 69.436 ;
        RECT 50.808 69.434 67.776 69.482 ;
        RECT 50.762 69.48 67.73 69.528 ;
        RECT 50.716 69.526 67.684 69.574 ;
        RECT 50.67 69.572 67.638 69.62 ;
        RECT 50.624 69.618 67.592 69.666 ;
        RECT 50.578 69.664 67.546 69.712 ;
        RECT 50.532 69.71 67.5 69.758 ;
        RECT 50.486 69.756 67.454 69.804 ;
        RECT 50.44 69.802 67.408 69.85 ;
        RECT 50.394 69.848 67.362 69.896 ;
        RECT 50.348 69.894 67.316 69.942 ;
        RECT 50.302 69.94 67.27 69.988 ;
        RECT 50.256 69.986 67.224 70.034 ;
        RECT 50.21 70.032 67.178 70.08 ;
        RECT 50.164 70.078 67.132 70.126 ;
        RECT 50.118 70.124 67.086 70.172 ;
        RECT 50.072 70.17 67.04 70.218 ;
        RECT 50.026 70.216 66.994 70.264 ;
        RECT 49.98 70.262 66.948 70.31 ;
        RECT 49.934 70.308 66.902 70.356 ;
        RECT 49.888 70.354 66.856 70.402 ;
        RECT 49.842 70.4 66.81 70.448 ;
        RECT 49.796 70.446 66.764 70.494 ;
        RECT 49.75 70.492 66.718 70.54 ;
        RECT 49.704 70.538 66.672 70.586 ;
        RECT 49.658 70.584 66.626 70.632 ;
        RECT 49.612 70.63 66.58 70.678 ;
        RECT 49.566 70.676 66.534 70.724 ;
        RECT 49.52 70.722 66.488 70.77 ;
        RECT 49.474 70.768 66.442 70.816 ;
        RECT 49.428 70.814 66.396 70.862 ;
        RECT 49.382 70.86 66.35 70.908 ;
        RECT 49.336 70.906 66.304 70.954 ;
        RECT 49.29 70.952 66.258 71 ;
        RECT 49.244 70.998 66.212 71.046 ;
        RECT 49.198 71.044 66.166 71.092 ;
        RECT 49.152 71.09 66.12 71.138 ;
        RECT 49.106 71.136 66.074 71.184 ;
        RECT 49.06 71.182 66.028 71.23 ;
        RECT 49.014 71.228 65.982 71.276 ;
        RECT 48.968 71.274 65.936 71.322 ;
        RECT 48.922 71.32 65.89 71.368 ;
        RECT 48.876 71.366 65.844 71.414 ;
        RECT 48.83 71.412 65.798 71.46 ;
        RECT 48.784 71.458 65.752 71.506 ;
        RECT 48.738 71.504 65.706 71.552 ;
        RECT 48.692 71.55 65.66 71.598 ;
        RECT 48.646 71.596 65.614 71.644 ;
        RECT 48.6 71.642 65.568 71.69 ;
        RECT 48.554 71.688 65.522 71.736 ;
        RECT 48.508 71.734 65.476 71.782 ;
        RECT 48.462 71.78 65.43 71.828 ;
        RECT 48.416 71.826 65.384 71.874 ;
        RECT 48.37 71.872 65.338 71.92 ;
        RECT 48.324 71.918 65.292 71.966 ;
        RECT 48.278 71.964 65.246 72.012 ;
        RECT 48.232 72.01 65.2 72.058 ;
        RECT 48.186 72.056 65.154 72.104 ;
        RECT 48.14 72.102 65.108 72.15 ;
        RECT 48.094 72.148 65.062 72.196 ;
        RECT 48.048 72.194 65.016 72.242 ;
        RECT 48.002 72.24 64.97 72.288 ;
        RECT 47.956 72.286 64.924 72.334 ;
        RECT 47.91 72.332 64.878 72.38 ;
        RECT 47.864 72.378 64.832 72.426 ;
        RECT 47.818 72.424 64.786 72.472 ;
        RECT 47.772 72.47 64.74 72.518 ;
        RECT 47.726 72.516 64.694 72.564 ;
        RECT 47.68 72.562 64.648 72.61 ;
        RECT 47.634 72.608 64.602 72.656 ;
        RECT 47.588 72.654 64.556 72.702 ;
        RECT 47.542 72.7 64.51 72.748 ;
        RECT 47.496 72.746 64.464 72.794 ;
        RECT 47.45 72.792 64.418 72.84 ;
        RECT 47.404 72.838 64.372 72.886 ;
        RECT 47.358 72.884 64.326 72.932 ;
        RECT 47.312 72.93 64.28 72.978 ;
        RECT 47.266 72.976 64.234 73.024 ;
        RECT 47.22 73.022 64.188 73.07 ;
        RECT 47.174 73.068 64.142 73.116 ;
        RECT 47.128 73.114 64.096 73.162 ;
        RECT 47.082 73.16 64.05 73.208 ;
        RECT 47.036 73.206 64.004 73.254 ;
        RECT 46.99 73.252 63.958 73.3 ;
        RECT 46.944 73.298 63.912 73.346 ;
        RECT 46.898 73.344 63.866 73.392 ;
        RECT 46.852 73.39 63.82 73.438 ;
        RECT 46.806 73.436 63.774 73.484 ;
        RECT 46.76 73.482 63.728 73.53 ;
        RECT 46.714 73.528 63.682 73.576 ;
        RECT 46.668 73.574 63.636 73.622 ;
        RECT 46.622 73.62 63.59 73.668 ;
        RECT 46.576 73.666 63.544 73.714 ;
        RECT 46.53 73.712 63.498 73.76 ;
        RECT 46.484 73.758 63.452 73.806 ;
        RECT 46.438 73.804 63.406 73.852 ;
        RECT 46.392 73.85 63.36 73.898 ;
        RECT 46.346 73.896 63.314 73.944 ;
        RECT 46.3 73.942 63.268 73.99 ;
        RECT 46.254 73.988 63.222 74.036 ;
        RECT 46.208 74.034 63.176 74.082 ;
        RECT 46.162 74.08 63.13 74.128 ;
        RECT 46.116 74.126 63.084 74.174 ;
        RECT 46.07 74.172 63.038 74.22 ;
        RECT 46.024 74.218 62.992 74.266 ;
        RECT 45.978 74.264 62.946 74.312 ;
        RECT 45.932 74.31 62.9 74.358 ;
        RECT 45.886 74.356 62.854 74.404 ;
        RECT 45.84 74.402 62.808 74.45 ;
        RECT 45.794 74.448 62.762 74.496 ;
        RECT 45.748 74.494 62.716 74.542 ;
        RECT 45.702 74.54 62.67 74.588 ;
        RECT 45.656 74.586 62.624 74.634 ;
        RECT 45.61 74.632 62.578 74.68 ;
        RECT 45.564 74.678 62.532 74.726 ;
        RECT 45.518 74.724 62.486 74.772 ;
        RECT 45.472 74.77 62.44 74.818 ;
        RECT 45.426 74.816 62.394 74.864 ;
        RECT 45.38 74.862 62.348 74.91 ;
        RECT 45.334 74.908 62.302 74.956 ;
        RECT 45.288 74.954 62.256 75.002 ;
        RECT 45.242 75 62.21 75.048 ;
        RECT 45.196 75.046 62.164 75.094 ;
        RECT 45.15 75.092 62.118 75.14 ;
        RECT 45.104 75.138 62.072 75.186 ;
        RECT 45.058 75.184 62.026 75.232 ;
        RECT 45.012 75.23 61.98 75.278 ;
        RECT 44.966 75.276 61.934 75.324 ;
        RECT 44.92 75.322 61.888 75.37 ;
        RECT 44.874 75.368 61.842 75.416 ;
        RECT 44.828 75.414 61.796 75.462 ;
        RECT 44.782 75.46 61.75 75.508 ;
        RECT 44.736 75.506 61.704 75.554 ;
        RECT 44.69 75.552 61.658 75.6 ;
        RECT 44.644 75.598 61.612 75.646 ;
        RECT 44.598 75.644 61.566 75.692 ;
        RECT 44.552 75.69 61.52 75.738 ;
        RECT 44.506 75.736 61.474 75.784 ;
        RECT 44.46 75.782 61.428 75.83 ;
        RECT 44.414 75.828 61.382 75.876 ;
        RECT 44.368 75.874 61.336 75.922 ;
        RECT 44.322 75.92 61.29 75.968 ;
        RECT 44.276 75.966 61.244 76.014 ;
        RECT 44.23 76.012 61.198 76.06 ;
        RECT 44.184 76.058 61.152 76.106 ;
        RECT 44.138 76.104 61.106 76.152 ;
        RECT 44.092 76.15 61.06 76.198 ;
        RECT 44.046 76.196 61.014 76.244 ;
        RECT 44 76.242 60.968 76.29 ;
        RECT 44 76.242 60.922 76.336 ;
        RECT 44 76.242 60.876 76.382 ;
        RECT 44 76.242 60.83 76.428 ;
        RECT 44 76.242 60.784 76.474 ;
        RECT 44 76.242 60.738 76.52 ;
        RECT 44 76.242 60.692 76.566 ;
        RECT 44 76.242 60.646 76.612 ;
        RECT 44 76.242 60.6 76.658 ;
        RECT 44 76.242 60.554 76.704 ;
        RECT 44 76.242 60.508 76.75 ;
        RECT 44 76.242 60.462 76.796 ;
        RECT 44 76.242 60.416 76.842 ;
        RECT 44 76.242 60.37 76.888 ;
        RECT 44 76.242 60.324 76.934 ;
        RECT 44 76.242 60.278 76.98 ;
        RECT 44 76.242 60.232 77.026 ;
        RECT 44 76.242 60.186 77.072 ;
        RECT 44 76.242 60.14 77.118 ;
        RECT 44 76.242 60.094 77.164 ;
        RECT 44 76.242 60.048 77.21 ;
        RECT 44 76.242 60.002 77.256 ;
        RECT 44 76.242 59.956 77.302 ;
        RECT 44 76.242 59.91 77.348 ;
        RECT 44 76.242 59.864 77.394 ;
        RECT 44 76.242 59.818 77.44 ;
        RECT 44 76.242 59.772 77.486 ;
        RECT 44 76.242 59.726 77.532 ;
        RECT 44 76.242 59.68 77.578 ;
        RECT 44 76.242 59.634 77.624 ;
        RECT 44 76.242 59.588 77.67 ;
        RECT 44 76.242 59.542 77.716 ;
        RECT 44 76.242 59.496 77.762 ;
        RECT 44 76.242 59.45 77.808 ;
        RECT 44 76.242 59.404 77.854 ;
        RECT 44 76.242 59.358 77.9 ;
        RECT 44 76.242 59.312 77.946 ;
        RECT 44 76.242 59.266 77.992 ;
        RECT 44 76.242 59.22 78.038 ;
        RECT 44 76.242 59.174 78.084 ;
        RECT 44 76.242 59.128 78.13 ;
        RECT 44 76.242 59.082 78.176 ;
        RECT 44 76.242 59.036 78.222 ;
        RECT 44 76.242 58.99 78.268 ;
        RECT 44 76.242 58.944 78.314 ;
        RECT 44 76.242 58.898 78.36 ;
        RECT 44 76.242 58.852 78.406 ;
        RECT 44 76.242 58.806 78.452 ;
        RECT 44 76.242 58.76 78.498 ;
        RECT 44 76.242 58.714 78.544 ;
        RECT 44 76.242 58.668 78.59 ;
        RECT 44 76.242 58.622 78.636 ;
        RECT 44 76.242 58.576 78.682 ;
        RECT 44 76.242 58.53 78.728 ;
        RECT 44 76.242 58.484 78.774 ;
        RECT 44 76.242 58.438 78.82 ;
        RECT 44 76.242 58.392 78.866 ;
        RECT 44 76.242 58.346 78.912 ;
        RECT 44 76.242 58.3 78.958 ;
        RECT 44 76.242 58.254 79.004 ;
        RECT 44 76.242 58.208 79.05 ;
        RECT 44 76.242 58.162 79.096 ;
        RECT 44 76.242 58.116 79.142 ;
        RECT 44 76.242 58.07 79.188 ;
        RECT 44 76.242 58.024 79.234 ;
        RECT 44 76.242 57.978 79.28 ;
        RECT 44 76.242 57.932 79.326 ;
        RECT 44 76.242 57.886 79.372 ;
        RECT 44 76.242 57.84 79.418 ;
        RECT 44 76.242 57.794 79.464 ;
        RECT 44 76.242 57.748 79.51 ;
        RECT 44 76.242 57.702 79.556 ;
        RECT 44 76.242 57.656 79.602 ;
        RECT 44 76.242 57.61 79.648 ;
        RECT 44 76.242 57.564 79.694 ;
        RECT 44 76.242 57.518 79.74 ;
        RECT 44 76.242 57.472 79.786 ;
        RECT 44 76.242 57.426 79.832 ;
        RECT 44 76.242 57.38 79.878 ;
        RECT 44 76.242 57.334 79.924 ;
        RECT 44 76.242 57.288 79.97 ;
        RECT 44 76.242 57.242 80.016 ;
        RECT 44 76.242 57.196 80.062 ;
        RECT 44 76.242 57.15 80.108 ;
        RECT 44 76.242 57.104 80.154 ;
        RECT 44 76.242 57.058 80.2 ;
        RECT 44 76.242 57.012 80.246 ;
        RECT 44 76.242 56.966 80.292 ;
        RECT 44 76.242 56.92 80.338 ;
        RECT 44 76.242 56.874 80.384 ;
        RECT 44 76.242 56.828 80.43 ;
        RECT 44 76.242 56.782 80.476 ;
        RECT 44 76.242 56.736 80.522 ;
        RECT 44 76.242 56.69 80.568 ;
        RECT 44 76.242 56.644 80.614 ;
        RECT 44 76.242 56.598 80.66 ;
        RECT 44 76.242 56.552 80.706 ;
        RECT 44 76.242 56.506 80.752 ;
        RECT 44 76.242 56.46 80.798 ;
        RECT 44 76.242 56.414 80.844 ;
        RECT 44 76.242 56.368 80.89 ;
        RECT 44 76.242 56.322 80.936 ;
        RECT 44 76.242 56.276 80.982 ;
        RECT 44 76.242 56.23 81.028 ;
        RECT 44 76.242 56.184 81.074 ;
        RECT 44 76.242 56.138 81.12 ;
        RECT 44 76.242 56.092 81.166 ;
        RECT 44 76.242 56.046 81.212 ;
        RECT 44 76.242 56 110 ;
        RECT 82.76 57.5 110 63.5 ;
        RECT 76.748 63.489 85.24 63.521 ;
        RECT 74.31 65.927 82.76 65.996 ;
        RECT 74.356 65.881 82.806 65.957 ;
        RECT 82.728 57.516 82.76 65.996 ;
        RECT 74.264 65.973 82.728 66.035 ;
        RECT 74.402 65.835 82.852 65.911 ;
        RECT 82.682 57.555 82.728 66.035 ;
        RECT 74.218 66.019 82.682 66.081 ;
        RECT 74.448 65.789 82.898 65.865 ;
        RECT 82.636 57.601 82.682 66.081 ;
        RECT 74.172 66.065 82.636 66.127 ;
        RECT 74.494 65.743 82.944 65.819 ;
        RECT 82.59 57.647 82.636 66.127 ;
        RECT 74.126 66.111 82.59 66.173 ;
        RECT 74.54 65.697 82.99 65.773 ;
        RECT 82.544 57.693 82.59 66.173 ;
        RECT 74.08 66.157 82.544 66.219 ;
        RECT 74.586 65.651 83.036 65.727 ;
        RECT 82.498 57.739 82.544 66.219 ;
        RECT 74.034 66.203 82.498 66.265 ;
        RECT 74.632 65.605 83.082 65.681 ;
        RECT 82.452 57.785 82.498 66.265 ;
        RECT 73.988 66.249 82.452 66.311 ;
        RECT 74.678 65.559 83.128 65.635 ;
        RECT 82.406 57.831 82.452 66.311 ;
        RECT 73.942 66.295 82.406 66.357 ;
        RECT 74.724 65.513 83.174 65.589 ;
        RECT 82.36 57.877 82.406 66.357 ;
        RECT 73.896 66.341 82.36 66.403 ;
        RECT 74.77 65.467 83.22 65.543 ;
        RECT 82.314 57.923 82.36 66.403 ;
        RECT 73.85 66.387 82.314 66.449 ;
        RECT 74.816 65.421 83.266 65.497 ;
        RECT 82.268 57.969 82.314 66.449 ;
        RECT 73.804 66.433 82.268 66.495 ;
        RECT 74.862 65.375 83.312 65.451 ;
        RECT 82.222 58.015 82.268 66.495 ;
        RECT 73.758 66.479 82.222 66.541 ;
        RECT 74.908 65.329 83.358 65.405 ;
        RECT 82.176 58.061 82.222 66.541 ;
        RECT 73.712 66.525 82.176 66.587 ;
        RECT 74.954 65.283 83.404 65.359 ;
        RECT 82.13 58.107 82.176 66.587 ;
        RECT 73.666 66.571 82.13 66.633 ;
        RECT 75 65.237 83.45 65.313 ;
        RECT 82.084 58.153 82.13 66.633 ;
        RECT 73.62 66.617 82.084 66.679 ;
        RECT 75.046 65.191 83.496 65.267 ;
        RECT 82.038 58.199 82.084 66.679 ;
        RECT 73.574 66.663 82.038 66.725 ;
        RECT 75.092 65.145 83.542 65.221 ;
        RECT 81.992 58.245 82.038 66.725 ;
        RECT 73.528 66.709 81.992 66.771 ;
        RECT 75.138 65.099 83.588 65.175 ;
        RECT 81.946 58.291 81.992 66.771 ;
        RECT 73.482 66.755 81.946 66.817 ;
        RECT 75.184 65.053 83.634 65.129 ;
        RECT 81.9 58.337 81.946 66.817 ;
        RECT 73.436 66.801 81.9 66.863 ;
        RECT 75.23 65.007 83.68 65.083 ;
        RECT 81.854 58.383 81.9 66.863 ;
        RECT 73.39 66.847 81.854 66.909 ;
        RECT 75.276 64.961 83.726 65.037 ;
        RECT 81.808 58.429 81.854 66.909 ;
        RECT 73.344 66.893 81.808 66.955 ;
        RECT 75.322 64.915 83.772 64.991 ;
        RECT 81.762 58.475 81.808 66.955 ;
        RECT 73.298 66.939 81.762 67.001 ;
        RECT 75.368 64.869 83.818 64.945 ;
        RECT 81.716 58.521 81.762 67.001 ;
        RECT 73.252 66.985 81.716 67.047 ;
        RECT 75.414 64.823 83.864 64.899 ;
        RECT 81.67 58.567 81.716 67.047 ;
        RECT 73.206 67.031 81.67 67.093 ;
        RECT 75.46 64.777 83.91 64.853 ;
        RECT 81.624 58.613 81.67 67.093 ;
        RECT 73.16 67.077 81.624 67.139 ;
        RECT 75.506 64.731 83.956 64.807 ;
        RECT 81.578 58.659 81.624 67.139 ;
        RECT 73.114 67.123 81.578 67.185 ;
        RECT 75.552 64.685 84.002 64.761 ;
        RECT 81.532 58.705 81.578 67.185 ;
        RECT 73.068 67.169 81.532 67.231 ;
        RECT 75.598 64.639 84.048 64.715 ;
        RECT 81.486 58.751 81.532 67.231 ;
        RECT 73.022 67.215 81.486 67.277 ;
        RECT 75.644 64.593 84.094 64.669 ;
        RECT 81.44 58.797 81.486 67.277 ;
        RECT 72.976 67.261 81.44 67.323 ;
        RECT 75.69 64.547 84.14 64.623 ;
        RECT 81.394 58.843 81.44 67.323 ;
        RECT 72.93 67.307 81.394 67.369 ;
        RECT 75.736 64.501 84.186 64.577 ;
        RECT 81.348 58.889 81.394 67.369 ;
        RECT 72.884 67.353 81.348 67.415 ;
        RECT 75.782 64.455 84.232 64.531 ;
        RECT 81.302 58.935 81.348 67.415 ;
        RECT 72.838 67.399 81.302 67.461 ;
        RECT 75.828 64.409 84.278 64.485 ;
        RECT 81.256 58.981 81.302 67.461 ;
        RECT 72.792 67.445 81.256 67.507 ;
        RECT 75.874 64.363 84.324 64.439 ;
        RECT 81.21 59.027 81.256 67.507 ;
        RECT 72.746 67.491 81.21 67.553 ;
        RECT 75.92 64.317 84.37 64.393 ;
        RECT 81.164 59.073 81.21 67.553 ;
        RECT 72.7 67.537 81.164 67.599 ;
        RECT 75.966 64.271 84.416 64.347 ;
        RECT 81.118 59.119 81.164 67.599 ;
        RECT 72.654 67.583 81.118 67.645 ;
        RECT 76.012 64.225 84.462 64.301 ;
        RECT 81.072 59.165 81.118 67.645 ;
        RECT 72.608 67.629 81.072 67.691 ;
        RECT 76.058 64.179 84.508 64.255 ;
        RECT 81.026 59.211 81.072 67.691 ;
        RECT 72.562 67.675 81.026 67.737 ;
        RECT 76.104 64.133 84.554 64.209 ;
        RECT 80.98 59.257 81.026 67.737 ;
        RECT 72.516 67.721 80.98 67.783 ;
        RECT 76.15 64.087 84.6 64.163 ;
        RECT 80.934 59.303 80.98 67.783 ;
        RECT 72.47 67.767 80.934 67.829 ;
        RECT 76.196 64.041 84.646 64.117 ;
        RECT 80.888 59.349 80.934 67.829 ;
        RECT 72.424 67.813 80.888 67.875 ;
        RECT 76.242 63.995 84.692 64.071 ;
        RECT 80.842 59.395 80.888 67.875 ;
        RECT 72.378 67.859 80.842 67.921 ;
        RECT 76.288 63.949 84.738 64.025 ;
        RECT 80.796 59.441 80.842 67.921 ;
        RECT 72.332 67.905 80.796 67.967 ;
        RECT 76.334 63.903 84.784 63.979 ;
        RECT 80.75 59.487 80.796 67.967 ;
        RECT 72.286 67.951 80.75 68.013 ;
        RECT 76.38 63.857 84.83 63.933 ;
        RECT 80.704 59.533 80.75 68.013 ;
        RECT 72.24 67.997 80.704 68.059 ;
        RECT 76.426 63.811 84.876 63.887 ;
        RECT 80.658 59.579 80.704 68.059 ;
        RECT 72.194 68.043 80.658 68.105 ;
        RECT 76.472 63.765 84.922 63.841 ;
        RECT 80.612 59.625 80.658 68.105 ;
        RECT 72.148 68.089 80.612 68.151 ;
        RECT 76.518 63.719 84.968 63.795 ;
        RECT 80.566 59.671 80.612 68.151 ;
        RECT 72.102 68.135 80.566 68.197 ;
        RECT 76.564 63.673 85.014 63.749 ;
        RECT 80.52 59.717 80.566 68.197 ;
        RECT 72.056 68.181 80.52 68.243 ;
        RECT 76.61 63.627 85.06 63.703 ;
        RECT 80.474 59.763 80.52 68.243 ;
        RECT 72.01 68.227 80.474 68.289 ;
        RECT 76.656 63.581 85.106 63.657 ;
        RECT 80.428 59.809 80.474 68.289 ;
        RECT 71.964 68.273 80.428 68.335 ;
        RECT 76.702 63.535 85.152 63.611 ;
        RECT 80.382 59.855 80.428 68.335 ;
        RECT 71.918 68.319 80.382 68.381 ;
        RECT 76.748 63.489 85.198 63.565 ;
        RECT 80.336 59.901 80.382 68.381 ;
        RECT 71.872 68.365 80.336 68.427 ;
        RECT 76.794 63.443 110 63.5 ;
        RECT 80.29 59.947 80.336 68.427 ;
        RECT 71.826 68.411 80.29 68.473 ;
        RECT 76.84 63.397 110 63.5 ;
        RECT 80.244 59.993 80.29 68.473 ;
        RECT 71.78 68.457 80.244 68.519 ;
        RECT 76.886 63.351 110 63.5 ;
        RECT 80.198 60.039 80.244 68.519 ;
        RECT 71.734 68.503 80.198 68.565 ;
        RECT 76.932 63.305 110 63.5 ;
        RECT 80.152 60.085 80.198 68.565 ;
        RECT 71.688 68.549 80.152 68.611 ;
        RECT 76.978 63.259 110 63.5 ;
        RECT 80.106 60.131 80.152 68.611 ;
        RECT 71.642 68.595 80.106 68.657 ;
        RECT 77.024 63.213 110 63.5 ;
        RECT 80.06 60.177 80.106 68.657 ;
        RECT 71.596 68.641 80.06 68.703 ;
        RECT 77.07 63.167 110 63.5 ;
        RECT 80.014 60.223 80.06 68.703 ;
        RECT 71.55 68.687 80.014 68.749 ;
        RECT 77.116 63.121 110 63.5 ;
        RECT 79.968 60.269 80.014 68.749 ;
        RECT 71.504 68.733 79.968 68.795 ;
        RECT 77.162 63.075 110 63.5 ;
        RECT 79.922 60.315 79.968 68.795 ;
        RECT 71.458 68.779 79.922 68.841 ;
        RECT 77.208 63.029 110 63.5 ;
        RECT 79.876 60.361 79.922 68.841 ;
        RECT 71.412 68.825 79.876 68.887 ;
        RECT 77.254 62.983 110 63.5 ;
        RECT 79.83 60.407 79.876 68.887 ;
        RECT 71.366 68.871 79.83 68.933 ;
        RECT 77.3 62.937 110 63.5 ;
        RECT 79.784 60.453 79.83 68.933 ;
        RECT 71.32 68.917 79.784 68.979 ;
        RECT 77.346 62.891 110 63.5 ;
        RECT 79.738 60.499 79.784 68.979 ;
        RECT 71.274 68.963 79.738 69.025 ;
        RECT 77.392 62.845 110 63.5 ;
        RECT 79.692 60.545 79.738 69.025 ;
        RECT 71.228 69.009 79.692 69.071 ;
        RECT 77.438 62.799 110 63.5 ;
        RECT 79.646 60.591 79.692 69.071 ;
        RECT 71.182 69.055 79.646 69.117 ;
        RECT 77.484 62.753 110 63.5 ;
        RECT 79.6 60.637 79.646 69.117 ;
        RECT 71.136 69.101 79.6 69.163 ;
        RECT 77.53 62.707 110 63.5 ;
        RECT 79.554 60.683 79.6 69.163 ;
        RECT 71.09 69.147 79.554 69.209 ;
        RECT 77.576 62.661 110 63.5 ;
        RECT 79.508 60.729 79.554 69.209 ;
        RECT 71.044 69.193 79.508 69.255 ;
        RECT 77.622 62.615 110 63.5 ;
        RECT 79.462 60.775 79.508 69.255 ;
        RECT 70.998 69.239 79.462 69.301 ;
        RECT 77.668 62.569 110 63.5 ;
        RECT 79.416 60.821 79.462 69.301 ;
        RECT 70.952 69.285 79.416 69.347 ;
        RECT 77.714 62.523 110 63.5 ;
        RECT 79.37 60.867 79.416 69.347 ;
        RECT 70.906 69.331 79.37 69.393 ;
        RECT 77.76 62.477 110 63.5 ;
        RECT 79.324 60.913 79.37 69.393 ;
        RECT 70.86 69.377 79.324 69.439 ;
        RECT 77.806 62.431 110 63.5 ;
        RECT 79.278 60.959 79.324 69.439 ;
        RECT 69.515 30.5 110 42.5 ;
        RECT 57.496 42.496 74.483 42.524 ;
        RECT 52.574 47.418 69.515 47.477 ;
        RECT 52.62 47.372 69.561 47.447 ;
        RECT 69.502 30.506 69.515 47.477 ;
        RECT 52.666 47.326 69.607 47.401 ;
        RECT 69.456 30.536 69.502 47.506 ;
        RECT 52.528 47.464 69.456 47.552 ;
        RECT 52.712 47.28 69.653 47.355 ;
        RECT 69.41 30.582 69.456 47.552 ;
        RECT 52.482 47.51 69.41 47.598 ;
        RECT 52.758 47.234 69.699 47.309 ;
        RECT 69.364 30.628 69.41 47.598 ;
        RECT 52.436 47.556 69.364 47.644 ;
        RECT 52.804 47.188 69.745 47.263 ;
        RECT 69.318 30.674 69.364 47.644 ;
        RECT 52.39 47.602 69.318 47.69 ;
        RECT 52.85 47.142 69.791 47.217 ;
        RECT 69.272 30.72 69.318 47.69 ;
        RECT 52.344 47.648 69.272 47.736 ;
        RECT 52.896 47.096 69.837 47.171 ;
        RECT 69.226 30.766 69.272 47.736 ;
        RECT 52.298 47.694 69.226 47.782 ;
        RECT 52.942 47.05 69.883 47.125 ;
        RECT 69.18 30.812 69.226 47.782 ;
        RECT 52.252 47.74 69.18 47.828 ;
        RECT 52.988 47.004 69.929 47.079 ;
        RECT 69.134 30.858 69.18 47.828 ;
        RECT 52.206 47.786 69.134 47.874 ;
        RECT 53.034 46.958 69.975 47.033 ;
        RECT 69.088 30.904 69.134 47.874 ;
        RECT 52.16 47.832 69.088 47.92 ;
        RECT 53.08 46.912 70.021 46.987 ;
        RECT 69.042 30.95 69.088 47.92 ;
        RECT 52.114 47.878 69.042 47.966 ;
        RECT 53.126 46.866 70.067 46.941 ;
        RECT 68.996 30.996 69.042 47.966 ;
        RECT 52.068 47.924 68.996 48.012 ;
        RECT 53.172 46.82 70.113 46.895 ;
        RECT 68.95 31.042 68.996 48.012 ;
        RECT 52.022 47.97 68.95 48.058 ;
        RECT 53.218 46.774 70.159 46.849 ;
        RECT 68.904 31.088 68.95 48.058 ;
        RECT 51.976 48.016 68.904 48.104 ;
        RECT 53.264 46.728 70.205 46.803 ;
        RECT 68.858 31.134 68.904 48.104 ;
        RECT 51.93 48.062 68.858 48.15 ;
        RECT 53.31 46.682 70.251 46.757 ;
        RECT 68.812 31.18 68.858 48.15 ;
        RECT 51.884 48.108 68.812 48.196 ;
        RECT 53.356 46.636 70.297 46.711 ;
        RECT 68.766 31.226 68.812 48.196 ;
        RECT 51.838 48.154 68.766 48.242 ;
        RECT 53.402 46.59 70.343 46.665 ;
        RECT 68.72 31.272 68.766 48.242 ;
        RECT 51.792 48.2 68.72 48.288 ;
        RECT 53.448 46.544 70.389 46.619 ;
        RECT 68.674 31.318 68.72 48.288 ;
        RECT 51.746 48.246 68.674 48.334 ;
        RECT 53.494 46.498 70.435 46.573 ;
        RECT 68.628 31.364 68.674 48.334 ;
        RECT 51.7 48.292 68.628 48.38 ;
        RECT 53.54 46.452 70.481 46.527 ;
        RECT 68.582 31.41 68.628 48.38 ;
        RECT 51.654 48.338 68.582 48.426 ;
        RECT 53.586 46.406 70.527 46.481 ;
        RECT 68.536 31.456 68.582 48.426 ;
        RECT 51.608 48.384 68.536 48.472 ;
        RECT 53.632 46.36 70.573 46.435 ;
        RECT 68.49 31.502 68.536 48.472 ;
        RECT 51.562 48.43 68.49 48.518 ;
        RECT 53.678 46.314 70.619 46.389 ;
        RECT 68.444 31.548 68.49 48.518 ;
        RECT 51.516 48.476 68.444 48.564 ;
        RECT 53.724 46.268 70.665 46.343 ;
        RECT 68.398 31.594 68.444 48.564 ;
        RECT 51.47 48.522 68.398 48.61 ;
        RECT 53.77 46.222 70.711 46.297 ;
        RECT 68.352 31.64 68.398 48.61 ;
        RECT 51.424 48.568 68.352 48.656 ;
        RECT 53.816 46.176 70.757 46.251 ;
        RECT 68.306 31.686 68.352 48.656 ;
        RECT 51.378 48.614 68.306 48.702 ;
        RECT 53.862 46.13 70.803 46.205 ;
        RECT 68.26 31.732 68.306 48.702 ;
        RECT 51.332 48.66 68.26 48.748 ;
        RECT 53.908 46.084 70.849 46.159 ;
        RECT 68.214 31.778 68.26 48.748 ;
        RECT 51.286 48.706 68.214 48.794 ;
        RECT 53.954 46.038 70.895 46.113 ;
        RECT 68.168 31.824 68.214 48.794 ;
        RECT 51.24 48.752 68.168 48.84 ;
        RECT 54 45.992 70.941 46.067 ;
        RECT 68.122 31.87 68.168 48.84 ;
        RECT 51.194 48.798 68.122 48.886 ;
        RECT 54.046 45.946 70.987 46.021 ;
        RECT 68.076 31.916 68.122 48.886 ;
        RECT 51.148 48.844 68.076 48.932 ;
        RECT 54.092 45.9 71.033 45.975 ;
        RECT 68.03 31.962 68.076 48.932 ;
        RECT 51.102 48.89 68.03 48.978 ;
        RECT 54.138 45.854 71.079 45.929 ;
        RECT 67.984 32.008 68.03 48.978 ;
        RECT 51.056 48.936 67.984 49.024 ;
        RECT 54.184 45.808 71.125 45.883 ;
        RECT 67.938 32.054 67.984 49.024 ;
        RECT 51.01 48.982 67.938 49.07 ;
        RECT 54.23 45.762 71.171 45.837 ;
        RECT 67.892 32.1 67.938 49.07 ;
        RECT 50.964 49.028 67.892 49.116 ;
        RECT 54.276 45.716 71.217 45.791 ;
        RECT 67.846 32.146 67.892 49.116 ;
        RECT 50.918 49.074 67.846 49.162 ;
        RECT 54.322 45.67 71.263 45.745 ;
        RECT 67.8 32.192 67.846 49.162 ;
        RECT 50.872 49.12 67.8 49.208 ;
        RECT 54.368 45.624 71.309 45.699 ;
        RECT 67.754 32.238 67.8 49.208 ;
        RECT 50.826 49.166 67.754 49.254 ;
        RECT 54.414 45.578 71.355 45.653 ;
        RECT 67.708 32.284 67.754 49.254 ;
        RECT 50.78 49.212 67.708 49.3 ;
        RECT 54.46 45.532 71.401 45.607 ;
        RECT 67.662 32.33 67.708 49.3 ;
        RECT 50.734 49.258 67.662 49.346 ;
        RECT 54.506 45.486 71.447 45.561 ;
        RECT 67.616 32.376 67.662 49.346 ;
        RECT 50.688 49.304 67.616 49.392 ;
        RECT 54.552 45.44 71.493 45.515 ;
        RECT 67.57 32.422 67.616 49.392 ;
        RECT 50.642 49.35 67.57 49.438 ;
        RECT 54.598 45.394 71.539 45.469 ;
        RECT 67.524 32.468 67.57 49.438 ;
        RECT 50.596 49.396 67.524 49.484 ;
        RECT 54.644 45.348 71.585 45.423 ;
        RECT 67.478 32.514 67.524 49.484 ;
        RECT 50.55 49.442 67.478 49.53 ;
        RECT 54.69 45.302 71.631 45.377 ;
        RECT 67.432 32.56 67.478 49.53 ;
        RECT 50.504 49.488 67.432 49.576 ;
        RECT 54.736 45.256 71.677 45.331 ;
        RECT 67.386 32.606 67.432 49.576 ;
        RECT 50.458 49.534 67.386 49.622 ;
        RECT 54.782 45.21 71.723 45.285 ;
        RECT 67.34 32.652 67.386 49.622 ;
        RECT 50.412 49.58 67.34 49.668 ;
        RECT 54.828 45.164 71.769 45.239 ;
        RECT 67.294 32.698 67.34 49.668 ;
        RECT 50.366 49.626 67.294 49.714 ;
        RECT 54.874 45.118 71.815 45.193 ;
        RECT 67.248 32.744 67.294 49.714 ;
        RECT 50.32 49.672 67.248 49.76 ;
        RECT 54.92 45.072 71.861 45.147 ;
        RECT 67.202 32.79 67.248 49.76 ;
        RECT 50.274 49.718 67.202 49.806 ;
        RECT 54.966 45.026 71.907 45.101 ;
        RECT 67.156 32.836 67.202 49.806 ;
        RECT 50.228 49.764 67.156 49.852 ;
        RECT 55.012 44.98 71.953 45.055 ;
        RECT 67.11 32.882 67.156 49.852 ;
        RECT 50.182 49.81 67.11 49.898 ;
        RECT 55.058 44.934 71.999 45.009 ;
        RECT 67.064 32.928 67.11 49.898 ;
        RECT 50.136 49.856 67.064 49.944 ;
        RECT 55.104 44.888 72.045 44.963 ;
        RECT 67.018 32.974 67.064 49.944 ;
        RECT 50.09 49.902 67.018 49.99 ;
        RECT 55.15 44.842 72.091 44.917 ;
        RECT 66.972 33.02 67.018 49.99 ;
        RECT 50.044 49.948 66.972 50.036 ;
        RECT 55.196 44.796 72.137 44.871 ;
        RECT 66.926 33.066 66.972 50.036 ;
        RECT 49.998 49.994 66.926 50.082 ;
        RECT 55.242 44.75 72.183 44.825 ;
        RECT 66.88 33.112 66.926 50.082 ;
        RECT 49.952 50.04 66.88 50.128 ;
        RECT 55.288 44.704 72.229 44.779 ;
        RECT 66.834 33.158 66.88 50.128 ;
        RECT 49.906 50.086 66.834 50.174 ;
        RECT 55.334 44.658 72.275 44.733 ;
        RECT 66.788 33.204 66.834 50.174 ;
        RECT 49.86 50.132 66.788 50.22 ;
        RECT 55.38 44.612 72.321 44.687 ;
        RECT 66.742 33.25 66.788 50.22 ;
        RECT 49.814 50.178 66.742 50.266 ;
        RECT 55.426 44.566 72.367 44.641 ;
        RECT 66.696 33.296 66.742 50.266 ;
        RECT 49.768 50.224 66.696 50.312 ;
        RECT 55.472 44.52 72.413 44.595 ;
        RECT 66.65 33.342 66.696 50.312 ;
        RECT 49.722 50.27 66.65 50.358 ;
        RECT 55.518 44.474 72.459 44.549 ;
        RECT 66.604 33.388 66.65 50.358 ;
        RECT 49.676 50.316 66.604 50.404 ;
        RECT 55.564 44.428 72.505 44.503 ;
        RECT 66.558 33.434 66.604 50.404 ;
        RECT 49.63 50.362 66.558 50.45 ;
        RECT 55.61 44.382 72.551 44.457 ;
        RECT 66.512 33.48 66.558 50.45 ;
        RECT 49.584 50.408 66.512 50.496 ;
        RECT 55.656 44.336 72.597 44.411 ;
        RECT 66.466 33.526 66.512 50.496 ;
        RECT 49.538 50.454 66.466 50.542 ;
        RECT 55.702 44.29 72.643 44.365 ;
        RECT 66.42 33.572 66.466 50.542 ;
        RECT 49.492 50.5 66.42 50.588 ;
        RECT 55.748 44.244 72.689 44.319 ;
        RECT 66.374 33.618 66.42 50.588 ;
        RECT 49.446 50.546 66.374 50.634 ;
        RECT 55.794 44.198 72.735 44.273 ;
        RECT 66.328 33.664 66.374 50.634 ;
        RECT 49.4 50.592 66.328 50.68 ;
        RECT 55.84 44.152 72.781 44.227 ;
        RECT 66.282 33.71 66.328 50.68 ;
        RECT 49.354 50.638 66.282 50.726 ;
        RECT 55.886 44.106 72.827 44.181 ;
        RECT 66.236 33.756 66.282 50.726 ;
        RECT 49.308 50.684 66.236 50.772 ;
        RECT 55.932 44.06 72.873 44.135 ;
        RECT 66.19 33.802 66.236 50.772 ;
        RECT 49.262 50.73 66.19 50.818 ;
        RECT 55.978 44.014 72.919 44.089 ;
        RECT 66.144 33.848 66.19 50.818 ;
        RECT 49.216 50.776 66.144 50.864 ;
        RECT 56.024 43.968 72.965 44.043 ;
        RECT 66.098 33.894 66.144 50.864 ;
        RECT 49.17 50.822 66.098 50.91 ;
        RECT 56.07 43.922 73.011 43.997 ;
        RECT 66.052 33.94 66.098 50.91 ;
        RECT 49.124 50.868 66.052 50.956 ;
        RECT 56.116 43.876 73.057 43.951 ;
        RECT 66.006 33.986 66.052 50.956 ;
        RECT 49.078 50.914 66.006 51.002 ;
        RECT 56.162 43.83 73.103 43.905 ;
        RECT 65.96 34.032 66.006 51.002 ;
        RECT 49.032 50.96 65.96 51.048 ;
        RECT 56.208 43.784 73.149 43.859 ;
        RECT 65.914 34.078 65.96 51.048 ;
        RECT 48.986 51.006 65.914 51.094 ;
        RECT 56.254 43.738 73.195 43.813 ;
        RECT 65.868 34.124 65.914 51.094 ;
        RECT 48.94 51.052 65.868 51.14 ;
        RECT 56.3 43.692 73.241 43.767 ;
        RECT 65.822 34.17 65.868 51.14 ;
        RECT 48.894 51.098 65.822 51.186 ;
        RECT 56.346 43.646 73.287 43.721 ;
        RECT 65.776 34.216 65.822 51.186 ;
        RECT 48.848 51.144 65.776 51.232 ;
        RECT 56.392 43.6 73.333 43.675 ;
        RECT 65.73 34.262 65.776 51.232 ;
        RECT 48.802 51.19 65.73 51.278 ;
        RECT 56.438 43.554 73.379 43.629 ;
        RECT 65.684 34.308 65.73 51.278 ;
        RECT 48.756 51.236 65.684 51.324 ;
        RECT 56.484 43.508 73.425 43.583 ;
        RECT 65.638 34.354 65.684 51.324 ;
        RECT 48.71 51.282 65.638 51.37 ;
        RECT 56.53 43.462 73.471 43.537 ;
        RECT 65.592 34.4 65.638 51.37 ;
        RECT 48.664 51.328 65.592 51.416 ;
        RECT 56.576 43.416 73.517 43.491 ;
        RECT 65.546 34.446 65.592 51.416 ;
        RECT 48.618 51.374 65.546 51.462 ;
        RECT 56.622 43.37 73.563 43.445 ;
        RECT 65.5 34.492 65.546 51.462 ;
        RECT 48.572 51.42 65.5 51.508 ;
        RECT 56.668 43.324 73.609 43.399 ;
        RECT 65.454 34.538 65.5 51.508 ;
        RECT 48.526 51.466 65.454 51.554 ;
        RECT 56.714 43.278 73.655 43.353 ;
        RECT 65.408 34.584 65.454 51.554 ;
        RECT 48.48 51.512 65.408 51.6 ;
        RECT 56.76 43.232 73.701 43.307 ;
        RECT 65.362 34.63 65.408 51.6 ;
        RECT 48.434 51.558 65.362 51.646 ;
        RECT 56.806 43.186 73.747 43.261 ;
        RECT 65.316 34.676 65.362 51.646 ;
        RECT 48.388 51.604 65.316 51.692 ;
        RECT 56.852 43.14 73.793 43.215 ;
        RECT 65.27 34.722 65.316 51.692 ;
        RECT 48.342 51.65 65.27 51.738 ;
        RECT 56.898 43.094 73.839 43.169 ;
        RECT 65.224 34.768 65.27 51.738 ;
        RECT 48.296 51.696 65.224 51.784 ;
        RECT 56.944 43.048 73.885 43.123 ;
        RECT 65.178 34.814 65.224 51.784 ;
        RECT 48.25 51.742 65.178 51.83 ;
        RECT 56.99 43.002 73.931 43.077 ;
        RECT 65.132 34.86 65.178 51.83 ;
        RECT 48.204 51.788 65.132 51.876 ;
        RECT 57.036 42.956 73.977 43.031 ;
        RECT 65.086 34.906 65.132 51.876 ;
        RECT 48.158 51.834 65.086 51.922 ;
        RECT 57.082 42.91 74.023 42.985 ;
        RECT 65.04 34.952 65.086 51.922 ;
        RECT 48.112 51.88 65.04 51.968 ;
        RECT 57.128 42.864 74.069 42.939 ;
        RECT 64.994 34.998 65.04 51.968 ;
        RECT 48.066 51.926 64.994 52.014 ;
        RECT 57.174 42.818 74.115 42.893 ;
        RECT 64.948 35.044 64.994 52.014 ;
        RECT 48.02 51.972 64.948 52.06 ;
        RECT 57.22 42.772 74.161 42.847 ;
        RECT 64.902 35.09 64.948 52.06 ;
        RECT 47.974 52.018 64.902 52.106 ;
        RECT 57.266 42.726 74.207 42.801 ;
        RECT 64.856 35.136 64.902 52.106 ;
        RECT 47.928 52.064 64.856 52.152 ;
        RECT 57.312 42.68 74.253 42.755 ;
        RECT 64.81 35.182 64.856 52.152 ;
        RECT 47.882 52.11 64.81 52.198 ;
        RECT 57.358 42.634 74.299 42.709 ;
        RECT 64.764 35.228 64.81 52.198 ;
        RECT 47.836 52.156 64.764 52.244 ;
        RECT 57.404 42.588 74.345 42.663 ;
        RECT 64.718 35.274 64.764 52.244 ;
        RECT 47.79 52.202 64.718 52.29 ;
        RECT 57.45 42.542 74.391 42.617 ;
        RECT 64.672 35.32 64.718 52.29 ;
        RECT 47.744 52.248 64.672 52.336 ;
        RECT 57.496 42.496 74.437 42.571 ;
        RECT 64.626 35.366 64.672 52.336 ;
        RECT 47.698 52.294 64.626 52.382 ;
        RECT 57.542 42.45 110 42.5 ;
        RECT 64.58 35.412 64.626 52.382 ;
        RECT 47.652 52.34 64.58 52.428 ;
        RECT 57.588 42.404 110 42.5 ;
        RECT 64.534 35.458 64.58 52.428 ;
        RECT 47.606 52.386 64.534 52.474 ;
        RECT 57.634 42.358 110 42.5 ;
        RECT 64.488 35.504 64.534 52.474 ;
        RECT 47.56 52.432 64.488 52.52 ;
        RECT 57.68 42.312 110 42.5 ;
        RECT 64.442 35.55 64.488 52.52 ;
        RECT 47.514 52.478 64.442 52.566 ;
        RECT 57.726 42.266 110 42.5 ;
        RECT 64.396 35.596 64.442 52.566 ;
        RECT 47.468 52.524 64.396 52.612 ;
        RECT 57.772 42.22 110 42.5 ;
        RECT 64.35 35.642 64.396 52.612 ;
        RECT 47.422 52.57 64.35 52.658 ;
        RECT 57.818 42.174 110 42.5 ;
        RECT 64.304 35.688 64.35 52.658 ;
        RECT 47.376 52.616 64.304 52.704 ;
        RECT 57.864 42.128 110 42.5 ;
        RECT 64.258 35.734 64.304 52.704 ;
        RECT 47.33 52.662 64.258 52.75 ;
        RECT 57.91 42.082 110 42.5 ;
        RECT 64.212 35.78 64.258 52.75 ;
        RECT 47.284 52.708 64.212 52.796 ;
        RECT 57.956 42.036 110 42.5 ;
        RECT 64.166 35.826 64.212 52.796 ;
        RECT 47.238 52.754 64.166 52.842 ;
        RECT 58.002 41.99 110 42.5 ;
        RECT 64.12 35.872 64.166 52.842 ;
        RECT 47.192 52.8 64.12 52.888 ;
        RECT 58.048 41.944 110 42.5 ;
        RECT 64.074 35.918 64.12 52.888 ;
        RECT 47.146 52.846 64.074 52.934 ;
        RECT 58.094 41.898 110 42.5 ;
        RECT 64.028 35.964 64.074 52.934 ;
        RECT 47.1 52.892 64.028 52.98 ;
        RECT 58.14 41.852 110 42.5 ;
        RECT 63.982 36.01 64.028 52.98 ;
        RECT 47.054 52.938 63.982 53.026 ;
        RECT 58.186 41.806 110 42.5 ;
        RECT 63.936 36.056 63.982 53.026 ;
        RECT 47.008 52.984 63.936 53.072 ;
        RECT 58.232 41.76 110 42.5 ;
        RECT 63.89 36.102 63.936 53.072 ;
        RECT 46.962 53.03 63.89 53.118 ;
        RECT 58.278 41.714 110 42.5 ;
        RECT 63.844 36.148 63.89 53.118 ;
        RECT 46.916 53.076 63.844 53.164 ;
        RECT 58.324 41.668 110 42.5 ;
        RECT 63.798 36.194 63.844 53.164 ;
        RECT 46.87 53.122 63.798 53.21 ;
        RECT 58.37 41.622 110 42.5 ;
        RECT 63.752 36.24 63.798 53.21 ;
        RECT 46.824 53.168 63.752 53.256 ;
        RECT 58.416 41.576 110 42.5 ;
        RECT 63.706 36.286 63.752 53.256 ;
        RECT 46.778 53.214 63.706 53.302 ;
        RECT 58.462 41.53 110 42.5 ;
        RECT 63.66 36.332 63.706 53.302 ;
        RECT 46.732 53.26 63.66 53.348 ;
        RECT 58.508 41.484 110 42.5 ;
        RECT 63.614 36.378 63.66 53.348 ;
        RECT 46.686 53.306 63.614 53.394 ;
        RECT 58.554 41.438 110 42.5 ;
        RECT 63.568 36.424 63.614 53.394 ;
        RECT 46.64 53.352 63.568 53.44 ;
        RECT 58.6 41.392 110 42.5 ;
        RECT 63.522 36.47 63.568 53.44 ;
        RECT 46.594 53.398 63.522 53.486 ;
        RECT 58.646 41.346 110 42.5 ;
        RECT 63.476 36.516 63.522 53.486 ;
        RECT 46.548 53.444 63.476 53.532 ;
        RECT 58.692 41.3 110 42.5 ;
        RECT 63.43 36.562 63.476 53.532 ;
        RECT 46.502 53.49 63.43 53.578 ;
        RECT 58.738 41.254 110 42.5 ;
        RECT 63.384 36.608 63.43 53.578 ;
        RECT 46.456 53.536 63.384 53.624 ;
        RECT 58.784 41.208 110 42.5 ;
        RECT 63.338 36.654 63.384 53.624 ;
        RECT 46.41 53.582 63.338 53.67 ;
        RECT 58.83 41.162 110 42.5 ;
        RECT 63.292 36.7 63.338 53.67 ;
        RECT 46.364 53.628 63.292 53.716 ;
        RECT 58.876 41.116 110 42.5 ;
        RECT 63.246 36.746 63.292 53.716 ;
        RECT 46.318 53.674 63.246 53.762 ;
        RECT 58.922 41.07 110 42.5 ;
        RECT 63.2 36.792 63.246 53.762 ;
        RECT 46.272 53.72 63.2 53.808 ;
        RECT 58.968 41.024 110 42.5 ;
        RECT 63.154 36.838 63.2 53.808 ;
        RECT 46.226 53.766 63.154 53.854 ;
        RECT 59.014 40.978 110 42.5 ;
        RECT 63.108 36.884 63.154 53.854 ;
        RECT 46.18 53.812 63.108 53.9 ;
        RECT 59.06 40.932 110 42.5 ;
        RECT 63.062 36.93 63.108 53.9 ;
        RECT 46.134 53.858 63.062 53.946 ;
        RECT 59.106 40.886 110 42.5 ;
        RECT 63.016 36.976 63.062 53.946 ;
        RECT 46.088 53.904 63.016 53.992 ;
        RECT 59.152 40.84 110 42.5 ;
        RECT 62.97 37.022 63.016 53.992 ;
        RECT 46.042 53.95 62.97 54.038 ;
        RECT 59.198 40.794 110 42.5 ;
        RECT 62.924 37.068 62.97 54.038 ;
        RECT 45.996 53.996 62.924 54.084 ;
        RECT 59.244 40.748 110 42.5 ;
        RECT 62.878 37.114 62.924 54.084 ;
        RECT 45.95 54.042 62.878 54.13 ;
        RECT 59.29 40.702 110 42.5 ;
        RECT 62.832 37.16 62.878 54.13 ;
        RECT 45.904 54.088 62.832 54.176 ;
        RECT 59.336 40.656 110 42.5 ;
        RECT 62.786 37.206 62.832 54.176 ;
        RECT 45.858 54.134 62.786 54.222 ;
        RECT 59.382 40.61 110 42.5 ;
        RECT 62.74 37.252 62.786 54.222 ;
        RECT 45.812 54.18 62.74 54.268 ;
        RECT 59.428 40.564 110 42.5 ;
        RECT 62.694 37.298 62.74 54.268 ;
        RECT 45.766 54.226 62.694 54.314 ;
        RECT 59.474 40.518 110 42.5 ;
        RECT 62.648 37.344 62.694 54.314 ;
        RECT 45.72 54.272 62.648 54.36 ;
        RECT 59.52 40.472 110 42.5 ;
        RECT 62.602 37.39 62.648 54.36 ;
        RECT 45.674 54.318 62.602 54.406 ;
        RECT 59.566 40.426 110 42.5 ;
        RECT 62.556 37.436 62.602 54.406 ;
        RECT 45.628 54.364 62.556 54.452 ;
        RECT 59.612 40.38 110 42.5 ;
        RECT 62.51 37.482 62.556 54.452 ;
        RECT 45.582 54.41 62.51 54.498 ;
        RECT 59.658 40.334 110 42.5 ;
        RECT 62.464 37.528 62.51 54.498 ;
        RECT 45.536 54.456 62.464 54.544 ;
        RECT 59.704 40.288 110 42.5 ;
        RECT 62.418 37.574 62.464 54.544 ;
        RECT 45.49 54.502 62.418 54.59 ;
        RECT 59.75 40.242 110 42.5 ;
        RECT 62.372 37.62 62.418 54.59 ;
        RECT 45.444 54.548 62.372 54.636 ;
        RECT 59.796 40.196 110 42.5 ;
        RECT 62.326 37.666 62.372 54.636 ;
        RECT 45.398 54.594 62.326 54.682 ;
        RECT 59.842 40.15 110 42.5 ;
        RECT 62.28 37.712 62.326 54.682 ;
        RECT 45.352 54.64 62.28 54.728 ;
        RECT 59.888 40.104 110 42.5 ;
        RECT 62.234 37.758 62.28 54.728 ;
        RECT 45.306 54.686 62.234 54.774 ;
        RECT 59.934 40.058 110 42.5 ;
        RECT 62.188 37.804 62.234 54.774 ;
        RECT 45.26 54.732 62.188 54.82 ;
        RECT 59.98 40.012 110 42.5 ;
        RECT 62.142 37.85 62.188 54.82 ;
        RECT 45.214 54.778 62.142 54.866 ;
        RECT 60.026 39.966 110 42.5 ;
        RECT 62.096 37.896 62.142 54.866 ;
        RECT 45.168 54.824 62.096 54.912 ;
        RECT 60.072 39.92 110 42.5 ;
        RECT 62.05 37.942 62.096 54.912 ;
        RECT 45.122 54.87 62.05 54.958 ;
        RECT 60.118 39.874 110 42.5 ;
        RECT 62.004 37.988 62.05 54.958 ;
        RECT 45.076 54.916 62.004 55.004 ;
        RECT 60.164 39.828 110 42.5 ;
        RECT 61.958 38.034 62.004 55.004 ;
        RECT 45.03 54.962 61.958 55.05 ;
        RECT 60.21 39.782 110 42.5 ;
        RECT 61.912 38.08 61.958 55.05 ;
        RECT 44.984 55.008 61.912 55.096 ;
        RECT 60.256 39.736 110 42.5 ;
        RECT 61.866 38.126 61.912 55.096 ;
        RECT 44.938 55.054 61.866 55.142 ;
        RECT 60.302 39.69 110 42.5 ;
        RECT 61.82 38.172 61.866 55.142 ;
        RECT 44.892 55.1 61.82 55.188 ;
        RECT 60.348 39.644 110 42.5 ;
        RECT 61.774 38.218 61.82 55.188 ;
        RECT 44.846 55.146 61.774 55.234 ;
        RECT 60.394 39.598 110 42.5 ;
        RECT 61.728 38.264 61.774 55.234 ;
        RECT 44.8 55.192 61.728 55.28 ;
        RECT 60.44 39.552 110 42.5 ;
        RECT 61.682 38.31 61.728 55.28 ;
        RECT 44.754 55.238 61.682 55.326 ;
        RECT 60.486 39.506 110 42.5 ;
        RECT 61.636 38.356 61.682 55.326 ;
        RECT 44.708 55.284 61.636 55.372 ;
        RECT 60.532 39.46 110 42.5 ;
        RECT 61.59 38.402 61.636 55.372 ;
        RECT 44.662 55.33 61.59 55.418 ;
        RECT 60.578 39.414 110 42.5 ;
        RECT 61.544 38.448 61.59 55.418 ;
        RECT 44.616 55.376 61.544 55.464 ;
        RECT 60.624 39.368 110 42.5 ;
        RECT 61.498 38.494 61.544 55.464 ;
        RECT 44.57 55.422 61.498 55.51 ;
        RECT 60.67 39.322 110 42.5 ;
        RECT 61.452 38.54 61.498 55.51 ;
        RECT 44.524 55.468 61.452 55.556 ;
        RECT 60.716 39.276 110 42.5 ;
        RECT 61.406 38.586 61.452 55.556 ;
        RECT 44.478 55.514 61.406 55.602 ;
        RECT 60.762 39.23 110 42.5 ;
        RECT 61.36 38.632 61.406 55.602 ;
        RECT 44.432 55.56 61.36 55.648 ;
        RECT 60.808 39.184 110 42.5 ;
        RECT 61.314 38.678 61.36 55.648 ;
        RECT 44.386 55.606 61.314 55.694 ;
        RECT 60.854 39.138 110 42.5 ;
        RECT 61.268 38.724 61.314 55.694 ;
        RECT 44.34 55.652 61.268 55.74 ;
        RECT 60.9 39.092 110 42.5 ;
        RECT 61.222 38.77 61.268 55.74 ;
        RECT 44.294 55.698 61.222 55.786 ;
        RECT 60.946 39.046 110 42.5 ;
        RECT 61.176 38.816 61.222 55.786 ;
        RECT 44.248 55.744 61.176 55.832 ;
        RECT 60.992 39 110 42.5 ;
        RECT 61.13 38.862 61.176 55.832 ;
        RECT 44.202 55.79 61.13 55.878 ;
        RECT 61.038 38.954 110 42.5 ;
        RECT 61.084 38.908 61.13 55.878 ;
        RECT 44.156 55.836 61.084 55.924 ;
        RECT 44.11 55.882 61.038 55.97 ;
        RECT 44.064 55.928 60.992 56.016 ;
        RECT 44.018 55.974 60.946 56.062 ;
        RECT 43.972 56.02 60.9 56.108 ;
        RECT 43.926 56.066 60.854 56.154 ;
        RECT 43.88 56.112 60.808 56.2 ;
        RECT 43.834 56.158 60.762 56.246 ;
        RECT 43.788 56.204 60.716 56.292 ;
        RECT 43.742 56.25 60.67 56.338 ;
        RECT 43.696 56.296 60.624 56.384 ;
        RECT 43.65 56.342 60.578 56.43 ;
        RECT 43.604 56.388 60.532 56.476 ;
        RECT 43.558 56.434 60.486 56.522 ;
        RECT 43.512 56.48 60.44 56.568 ;
        RECT 43.466 56.526 60.394 56.614 ;
        RECT 43.42 56.572 60.348 56.66 ;
        RECT 43.374 56.618 60.302 56.706 ;
        RECT 43.328 56.664 60.256 56.752 ;
        RECT 43.282 56.71 60.21 56.798 ;
        RECT 43.236 56.756 60.164 56.844 ;
        RECT 43.19 56.802 60.118 56.89 ;
        RECT 43.144 56.848 60.072 56.936 ;
        RECT 43.098 56.894 60.026 56.982 ;
        RECT 43.052 56.94 59.98 57.028 ;
        RECT 43.006 56.986 59.934 57.074 ;
        RECT 42.96 57.032 59.888 57.12 ;
        RECT 42.914 57.078 59.842 57.166 ;
        RECT 42.868 57.124 59.796 57.212 ;
        RECT 42.822 57.17 59.75 57.258 ;
        RECT 42.776 57.216 59.704 57.304 ;
        RECT 42.73 57.262 59.658 57.35 ;
        RECT 42.684 57.308 59.612 57.396 ;
        RECT 42.638 57.354 59.566 57.442 ;
        RECT 42.592 57.4 59.52 57.488 ;
        RECT 42.5 57.492 59.474 57.534 ;
        RECT 42.546 57.446 59.474 57.534 ;
        RECT 42.46 57.535 59.428 57.58 ;
        RECT 42.414 57.578 59.382 57.626 ;
        RECT 42.368 57.624 59.336 57.672 ;
        RECT 42.322 57.67 59.29 57.718 ;
        RECT 42.276 57.716 59.244 57.764 ;
        RECT 42.23 57.762 59.198 57.81 ;
        RECT 42.184 57.808 59.152 57.856 ;
        RECT 42.138 57.854 59.106 57.902 ;
        RECT 42.092 57.9 59.06 57.948 ;
        RECT 42.046 57.946 59.014 57.994 ;
        RECT 42 57.992 58.968 58.04 ;
        RECT 41.954 58.038 58.922 58.086 ;
        RECT 41.908 58.084 58.876 58.132 ;
        RECT 41.862 58.13 58.83 58.178 ;
        RECT 41.816 58.176 58.784 58.224 ;
        RECT 41.77 58.222 58.738 58.27 ;
        RECT 41.724 58.268 58.692 58.316 ;
        RECT 41.678 58.314 58.646 58.362 ;
        RECT 41.632 58.36 58.6 58.408 ;
        RECT 41.586 58.406 58.554 58.454 ;
        RECT 41.54 58.452 58.508 58.5 ;
        RECT 41.494 58.498 58.462 58.546 ;
        RECT 41.448 58.544 58.416 58.592 ;
        RECT 41.402 58.59 58.37 58.638 ;
        RECT 41.356 58.636 58.324 58.684 ;
        RECT 41.31 58.682 58.278 58.73 ;
        RECT 41.264 58.728 58.232 58.776 ;
        RECT 41.218 58.774 58.186 58.822 ;
        RECT 41.172 58.82 58.14 58.868 ;
        RECT 41.126 58.866 58.094 58.914 ;
        RECT 41.08 58.912 58.048 58.96 ;
        RECT 41.034 58.958 58.002 59.006 ;
        RECT 40.988 59.004 57.956 59.052 ;
        RECT 40.942 59.05 57.91 59.098 ;
        RECT 40.896 59.096 57.864 59.144 ;
        RECT 40.85 59.142 57.818 59.19 ;
        RECT 40.804 59.188 57.772 59.236 ;
        RECT 40.758 59.234 57.726 59.282 ;
        RECT 40.712 59.28 57.68 59.328 ;
        RECT 40.666 59.326 57.634 59.374 ;
        RECT 40.62 59.372 57.588 59.42 ;
        RECT 40.574 59.418 57.542 59.466 ;
        RECT 40.528 59.464 57.496 59.512 ;
        RECT 40.482 59.51 57.45 59.558 ;
        RECT 40.436 59.556 57.404 59.604 ;
        RECT 40.39 59.602 57.358 59.65 ;
        RECT 40.344 59.648 57.312 59.696 ;
        RECT 40.298 59.694 57.266 59.742 ;
        RECT 40.252 59.74 57.22 59.788 ;
        RECT 40.206 59.786 57.174 59.834 ;
        RECT 40.16 59.832 57.128 59.88 ;
        RECT 40.114 59.878 57.082 59.926 ;
        RECT 40.068 59.924 57.036 59.972 ;
        RECT 40.022 59.97 56.99 60.018 ;
        RECT 39.976 60.016 56.944 60.064 ;
        RECT 39.93 60.062 56.898 60.11 ;
        RECT 39.884 60.108 56.852 60.156 ;
        RECT 39.838 60.154 56.806 60.202 ;
        RECT 39.792 60.2 56.76 60.248 ;
        RECT 39.746 60.246 56.714 60.294 ;
        RECT 39.7 60.292 56.668 60.34 ;
        RECT 39.654 60.338 56.622 60.386 ;
        RECT 39.608 60.384 56.576 60.432 ;
        RECT 39.562 60.43 56.53 60.478 ;
        RECT 39.516 60.476 56.484 60.524 ;
        RECT 39.47 60.522 56.438 60.57 ;
        RECT 39.424 60.568 56.392 60.616 ;
        RECT 39.378 60.614 56.346 60.662 ;
        RECT 39.332 60.66 56.3 60.708 ;
        RECT 39.286 60.706 56.254 60.754 ;
        RECT 39.24 60.752 56.208 60.8 ;
        RECT 39.194 60.798 56.162 60.846 ;
        RECT 39.148 60.844 56.116 60.892 ;
        RECT 39.102 60.89 56.07 60.938 ;
        RECT 39.056 60.936 56.024 60.984 ;
        RECT 39.01 60.982 55.978 61.03 ;
        RECT 38.964 61.028 55.932 61.076 ;
        RECT 38.918 61.074 55.886 61.122 ;
        RECT 38.872 61.12 55.84 61.168 ;
        RECT 38.826 61.166 55.794 61.214 ;
        RECT 38.78 61.212 55.748 61.26 ;
        RECT 38.734 61.258 55.702 61.306 ;
        RECT 38.688 61.304 55.656 61.352 ;
        RECT 38.642 61.35 55.61 61.398 ;
        RECT 38.596 61.396 55.564 61.444 ;
        RECT 38.55 61.442 55.518 61.49 ;
        RECT 38.504 61.488 55.472 61.536 ;
        RECT 38.458 61.534 55.426 61.582 ;
        RECT 38.412 61.58 55.38 61.628 ;
        RECT 38.366 61.626 55.334 61.674 ;
        RECT 38.32 61.672 55.288 61.72 ;
        RECT 38.274 61.718 55.242 61.766 ;
        RECT 38.228 61.764 55.196 61.812 ;
        RECT 38.182 61.81 55.15 61.858 ;
        RECT 38.136 61.856 55.104 61.904 ;
        RECT 38.09 61.902 55.058 61.95 ;
        RECT 38.044 61.948 55.012 61.996 ;
        RECT 37.998 61.994 54.966 62.042 ;
        RECT 37.952 62.04 54.92 62.088 ;
        RECT 37.906 62.086 54.874 62.134 ;
        RECT 37.86 62.132 54.828 62.18 ;
        RECT 37.814 62.178 54.782 62.226 ;
        RECT 37.768 62.224 54.736 62.272 ;
        RECT 37.722 62.27 54.69 62.318 ;
        RECT 37.676 62.316 54.644 62.364 ;
        RECT 37.63 62.362 54.598 62.41 ;
        RECT 37.584 62.408 54.552 62.456 ;
        RECT 37.538 62.454 54.506 62.502 ;
        RECT 37.492 62.5 54.46 62.548 ;
        RECT 37.446 62.546 54.414 62.594 ;
        RECT 37.4 62.592 54.368 62.64 ;
        RECT 37.354 62.638 54.322 62.686 ;
        RECT 37.308 62.684 54.276 62.732 ;
        RECT 37.262 62.73 54.23 62.778 ;
        RECT 37.216 62.776 54.184 62.824 ;
        RECT 37.17 62.822 54.138 62.87 ;
        RECT 37.124 62.868 54.092 62.916 ;
        RECT 37.078 62.914 54.046 62.962 ;
        RECT 37.032 62.96 54 63.008 ;
        RECT 36.986 63.006 53.954 63.054 ;
        RECT 36.94 63.052 53.908 63.1 ;
        RECT 36.894 63.098 53.862 63.146 ;
        RECT 36.848 63.144 53.816 63.192 ;
        RECT 36.802 63.19 53.77 63.238 ;
        RECT 36.756 63.236 53.724 63.284 ;
        RECT 36.71 63.282 53.678 63.33 ;
        RECT 36.664 63.328 53.632 63.376 ;
        RECT 36.618 63.374 53.586 63.422 ;
        RECT 36.572 63.42 53.54 63.468 ;
        RECT 36.526 63.466 53.494 63.514 ;
        RECT 36.48 63.512 53.448 63.56 ;
        RECT 36.434 63.558 53.402 63.606 ;
        RECT 36.388 63.604 53.356 63.652 ;
        RECT 36.342 63.65 53.31 63.698 ;
        RECT 36.296 63.696 53.264 63.744 ;
        RECT 36.25 63.742 53.218 63.79 ;
        RECT 36.204 63.788 53.172 63.836 ;
        RECT 36.158 63.834 53.126 63.882 ;
        RECT 36.112 63.88 53.08 63.928 ;
        RECT 36.066 63.926 53.034 63.974 ;
        RECT 36.02 63.972 52.988 64.02 ;
        RECT 35.974 64.018 52.942 64.066 ;
        RECT 35.928 64.064 52.896 64.112 ;
        RECT 35.882 64.11 52.85 64.158 ;
        RECT 35.836 64.156 52.804 64.204 ;
        RECT 35.79 64.202 52.758 64.25 ;
        RECT 35.744 64.248 52.712 64.296 ;
        RECT 35.698 64.294 52.666 64.342 ;
        RECT 35.652 64.34 52.62 64.388 ;
        RECT 35.606 64.386 52.574 64.434 ;
        RECT 35.56 64.432 52.528 64.48 ;
        RECT 35.514 64.478 52.482 64.526 ;
        RECT 35.468 64.524 52.436 64.572 ;
        RECT 35.422 64.57 52.39 64.618 ;
        RECT 35.376 64.616 52.344 64.664 ;
        RECT 35.33 64.662 52.298 64.71 ;
        RECT 35.284 64.708 52.252 64.756 ;
        RECT 35.238 64.754 52.206 64.802 ;
        RECT 35.192 64.8 52.16 64.848 ;
        RECT 35.146 64.846 52.114 64.894 ;
        RECT 35.1 64.892 52.068 64.94 ;
        RECT 35.054 64.938 52.022 64.986 ;
        RECT 35.008 64.984 51.976 65.032 ;
        RECT 34.962 65.03 51.93 65.078 ;
        RECT 34.916 65.076 51.884 65.124 ;
        RECT 34.87 65.122 51.838 65.17 ;
        RECT 34.824 65.168 51.792 65.216 ;
        RECT 34.778 65.214 51.746 65.262 ;
        RECT 34.732 65.26 51.7 65.308 ;
        RECT 34.686 65.306 51.654 65.354 ;
        RECT 34.64 65.352 51.608 65.4 ;
        RECT 34.594 65.398 51.562 65.446 ;
        RECT 34.548 65.444 51.516 65.492 ;
        RECT 34.502 65.49 51.47 65.538 ;
        RECT 34.456 65.536 51.424 65.584 ;
        RECT 34.41 65.582 51.378 65.63 ;
        RECT 34.364 65.628 51.332 65.676 ;
        RECT 34.318 65.674 51.286 65.722 ;
        RECT 34.272 65.72 51.24 65.768 ;
        RECT 34.226 65.766 51.194 65.814 ;
        RECT 34.18 65.812 51.148 65.86 ;
        RECT 34.134 65.858 51.102 65.906 ;
        RECT 34.088 65.904 51.056 65.952 ;
        RECT 34.042 65.95 51.01 65.998 ;
        RECT 33.996 65.996 50.964 66.044 ;
        RECT 33.95 66.042 50.918 66.09 ;
        RECT 33.904 66.088 50.872 66.136 ;
        RECT 33.858 66.134 50.826 66.182 ;
        RECT 33.812 66.18 50.78 66.228 ;
        RECT 33.766 66.226 50.734 66.274 ;
        RECT 33.72 66.272 50.688 66.32 ;
        RECT 33.674 66.318 50.642 66.366 ;
        RECT 33.628 66.364 50.596 66.412 ;
        RECT 33.582 66.41 50.55 66.458 ;
        RECT 33.536 66.456 50.504 66.504 ;
        RECT 33.49 66.502 50.458 66.55 ;
        RECT 33.444 66.548 50.412 66.596 ;
        RECT 33.398 66.594 50.366 66.642 ;
        RECT 33.352 66.64 50.32 66.688 ;
        RECT 33.306 66.686 50.274 66.734 ;
        RECT 33.26 66.732 50.228 66.78 ;
        RECT 33.214 66.778 50.182 66.826 ;
        RECT 33.168 66.824 50.136 66.872 ;
        RECT 33.122 66.87 50.09 66.918 ;
        RECT 33.076 66.916 50.044 66.964 ;
        RECT 33.03 66.962 49.998 67.01 ;
        RECT 32.984 67.008 49.952 67.056 ;
        RECT 32.938 67.054 49.906 67.102 ;
        RECT 32.892 67.1 49.86 67.148 ;
        RECT 32.846 67.146 49.814 67.194 ;
        RECT 32.8 67.192 49.768 67.24 ;
        RECT 32.754 67.238 49.722 67.286 ;
        RECT 32.708 67.284 49.676 67.332 ;
        RECT 32.662 67.33 49.63 67.378 ;
        RECT 32.616 67.376 49.584 67.424 ;
        RECT 32.57 67.422 49.538 67.47 ;
        RECT 32.524 67.468 49.492 67.516 ;
        RECT 32.478 67.514 49.446 67.562 ;
        RECT 32.432 67.56 49.4 67.608 ;
        RECT 32.386 67.606 49.354 67.654 ;
        RECT 32.34 67.652 49.308 67.7 ;
        RECT 32.294 67.698 49.262 67.746 ;
        RECT 32.248 67.744 49.216 67.792 ;
        RECT 32.202 67.79 49.17 67.838 ;
        RECT 32.156 67.836 49.124 67.884 ;
        RECT 32.11 67.882 49.078 67.93 ;
        RECT 32.064 67.928 49.032 67.976 ;
        RECT 32.018 67.974 48.986 68.022 ;
        RECT 31.972 68.02 48.94 68.068 ;
        RECT 31.926 68.066 48.894 68.114 ;
        RECT 31.88 68.112 48.848 68.16 ;
        RECT 31.834 68.158 48.802 68.206 ;
        RECT 31.788 68.204 48.756 68.252 ;
        RECT 31.742 68.25 48.71 68.298 ;
        RECT 31.696 68.296 48.664 68.344 ;
        RECT 31.65 68.342 48.618 68.39 ;
        RECT 31.604 68.388 48.572 68.436 ;
        RECT 31.558 68.434 48.526 68.482 ;
        RECT 31.512 68.48 48.48 68.528 ;
        RECT 31.466 68.526 48.434 68.574 ;
        RECT 31.42 68.572 48.388 68.62 ;
        RECT 31.374 68.618 48.342 68.666 ;
        RECT 31.328 68.664 48.296 68.712 ;
        RECT 31.282 68.71 48.25 68.758 ;
        RECT 31.236 68.756 48.204 68.804 ;
        RECT 31.19 68.802 48.158 68.85 ;
        RECT 31.144 68.848 48.112 68.896 ;
        RECT 31.098 68.894 48.066 68.942 ;
        RECT 31.052 68.94 48.02 68.988 ;
        RECT 31.006 68.986 47.974 69.034 ;
        RECT 30.96 69.032 47.928 69.08 ;
        RECT 30.914 69.078 47.882 69.126 ;
        RECT 30.868 69.124 47.836 69.172 ;
        RECT 30.822 69.17 47.79 69.218 ;
        RECT 30.776 69.216 47.744 69.264 ;
        RECT 30.73 69.262 47.698 69.31 ;
        RECT 30.684 69.308 47.652 69.356 ;
        RECT 30.638 69.354 47.606 69.402 ;
        RECT 30.592 69.4 47.56 69.448 ;
        RECT 30.546 69.446 47.514 69.494 ;
        RECT 30.5 69.492 47.468 69.54 ;
        RECT 30.5 69.492 47.422 69.586 ;
        RECT 30.5 69.492 47.376 69.632 ;
        RECT 30.5 69.492 47.33 69.678 ;
        RECT 30.5 69.492 47.284 69.724 ;
        RECT 30.5 69.492 47.238 69.77 ;
        RECT 30.5 69.492 47.192 69.816 ;
        RECT 30.5 69.492 47.146 69.862 ;
        RECT 30.5 69.492 47.1 69.908 ;
        RECT 30.5 69.492 47.054 69.954 ;
        RECT 30.5 69.492 47.008 70 ;
        RECT 30.5 69.492 46.962 70.046 ;
        RECT 30.5 69.492 46.916 70.092 ;
        RECT 30.5 69.492 46.87 70.138 ;
        RECT 30.5 69.492 46.824 70.184 ;
        RECT 30.5 69.492 46.778 70.23 ;
        RECT 30.5 69.492 46.732 70.276 ;
        RECT 30.5 69.492 46.686 70.322 ;
        RECT 30.5 69.492 46.64 70.368 ;
        RECT 30.5 69.492 46.594 70.414 ;
        RECT 30.5 69.492 46.548 70.46 ;
        RECT 30.5 69.492 46.502 70.506 ;
        RECT 30.5 69.492 46.456 70.552 ;
        RECT 30.5 69.492 46.41 70.598 ;
        RECT 30.5 69.492 46.364 70.644 ;
        RECT 30.5 69.492 46.318 70.69 ;
        RECT 30.5 69.492 46.272 70.736 ;
        RECT 30.5 69.492 46.226 70.782 ;
        RECT 30.5 69.492 46.18 70.828 ;
        RECT 30.5 69.492 46.134 70.874 ;
        RECT 30.5 69.492 46.088 70.92 ;
        RECT 30.5 69.492 46.042 70.966 ;
        RECT 30.5 69.492 45.996 71.012 ;
        RECT 30.5 69.492 45.95 71.058 ;
        RECT 30.5 69.492 45.904 71.104 ;
        RECT 30.5 69.492 45.858 71.15 ;
        RECT 30.5 69.492 45.812 71.196 ;
        RECT 30.5 69.492 45.766 71.242 ;
        RECT 30.5 69.492 45.72 71.288 ;
        RECT 30.5 69.492 45.674 71.334 ;
        RECT 30.5 69.492 45.628 71.38 ;
        RECT 30.5 69.492 45.582 71.426 ;
        RECT 30.5 69.492 45.536 71.472 ;
        RECT 30.5 69.492 45.49 71.518 ;
        RECT 30.5 69.492 45.444 71.564 ;
        RECT 30.5 69.492 45.398 71.61 ;
        RECT 30.5 69.492 45.352 71.656 ;
        RECT 30.5 69.492 45.306 71.702 ;
        RECT 30.5 69.492 45.26 71.748 ;
        RECT 30.5 69.492 45.214 71.794 ;
        RECT 30.5 69.492 45.168 71.84 ;
        RECT 30.5 69.492 45.122 71.886 ;
        RECT 30.5 69.492 45.076 71.932 ;
        RECT 30.5 69.492 45.03 71.978 ;
        RECT 30.5 69.492 44.984 72.024 ;
        RECT 30.5 69.492 44.938 72.07 ;
        RECT 30.5 69.492 44.892 72.116 ;
        RECT 30.5 69.492 44.846 72.162 ;
        RECT 30.5 69.492 44.8 72.208 ;
        RECT 30.5 69.492 44.754 72.254 ;
        RECT 30.5 69.492 44.708 72.3 ;
        RECT 30.5 69.492 44.662 72.346 ;
        RECT 30.5 69.492 44.616 72.392 ;
        RECT 30.5 69.492 44.57 72.438 ;
        RECT 30.5 69.492 44.524 72.484 ;
        RECT 30.5 69.492 44.478 72.53 ;
        RECT 30.5 69.492 44.432 72.576 ;
        RECT 30.5 69.492 44.386 72.622 ;
        RECT 30.5 69.492 44.34 72.668 ;
        RECT 30.5 69.492 44.294 72.714 ;
        RECT 30.5 69.492 44.248 72.76 ;
        RECT 30.5 69.492 44.202 72.806 ;
        RECT 30.5 69.492 44.156 72.852 ;
        RECT 30.5 69.492 44.11 72.898 ;
        RECT 30.5 69.492 44.064 72.944 ;
        RECT 30.5 69.492 44.018 72.99 ;
        RECT 30.5 69.492 43.972 73.036 ;
        RECT 30.5 69.492 43.926 73.082 ;
        RECT 30.5 69.492 43.88 73.128 ;
        RECT 30.5 69.492 43.834 73.174 ;
        RECT 30.5 69.492 43.788 73.22 ;
        RECT 30.5 69.492 43.742 73.266 ;
        RECT 30.5 69.492 43.696 73.312 ;
        RECT 30.5 69.492 43.65 73.358 ;
        RECT 30.5 69.492 43.604 73.404 ;
        RECT 30.5 69.492 43.558 73.45 ;
        RECT 30.5 69.492 43.512 73.496 ;
        RECT 30.5 69.492 43.466 73.542 ;
        RECT 30.5 69.492 43.42 73.588 ;
        RECT 30.5 69.492 43.374 73.634 ;
        RECT 30.5 69.492 43.328 73.68 ;
        RECT 30.5 69.492 43.282 73.726 ;
        RECT 30.5 69.492 43.236 73.772 ;
        RECT 30.5 69.492 43.19 73.818 ;
        RECT 30.5 69.492 43.144 73.864 ;
        RECT 30.5 69.492 43.098 73.91 ;
        RECT 30.5 69.492 43.052 73.956 ;
        RECT 30.5 69.492 43.006 74.002 ;
        RECT 30.5 69.492 42.96 74.048 ;
        RECT 30.5 69.492 42.914 74.094 ;
        RECT 30.5 69.492 42.868 74.14 ;
        RECT 30.5 69.492 42.822 74.186 ;
        RECT 30.5 69.492 42.776 74.232 ;
        RECT 30.5 69.492 42.73 74.278 ;
        RECT 30.5 69.492 42.684 74.324 ;
        RECT 30.5 69.492 42.638 74.37 ;
        RECT 30.5 69.492 42.592 74.416 ;
        RECT 30.5 69.492 42.546 74.462 ;
        RECT 30.5 69.492 42.5 110 ;
        RECT 76.265 44 110 56 ;
        RECT 59.312 60.93 76.265 60.983 ;
        RECT 59.358 60.884 76.311 60.947 ;
        RECT 76.24 44.012 76.265 60.983 ;
        RECT 59.404 60.838 76.357 60.901 ;
        RECT 76.194 44.048 76.24 61.018 ;
        RECT 59.266 60.976 76.194 61.064 ;
        RECT 59.45 60.792 76.403 60.855 ;
        RECT 76.148 44.094 76.194 61.064 ;
        RECT 59.22 61.022 76.148 61.11 ;
        RECT 59.496 60.746 76.449 60.809 ;
        RECT 76.102 44.14 76.148 61.11 ;
        RECT 59.174 61.068 76.102 61.156 ;
        RECT 59.542 60.7 76.495 60.763 ;
        RECT 76.056 44.186 76.102 61.156 ;
        RECT 59.128 61.114 76.056 61.202 ;
        RECT 59.588 60.654 76.541 60.717 ;
        RECT 76.01 44.232 76.056 61.202 ;
        RECT 59.082 61.16 76.01 61.248 ;
        RECT 59.634 60.608 76.587 60.671 ;
        RECT 75.964 44.278 76.01 61.248 ;
        RECT 59.036 61.206 75.964 61.294 ;
        RECT 59.68 60.562 76.633 60.625 ;
        RECT 75.918 44.324 75.964 61.294 ;
        RECT 58.99 61.252 75.918 61.34 ;
        RECT 59.726 60.516 76.679 60.579 ;
        RECT 75.872 44.37 75.918 61.34 ;
        RECT 58.944 61.298 75.872 61.386 ;
        RECT 59.772 60.47 76.725 60.533 ;
        RECT 75.826 44.416 75.872 61.386 ;
        RECT 58.898 61.344 75.826 61.432 ;
        RECT 59.818 60.424 76.771 60.487 ;
        RECT 75.78 44.462 75.826 61.432 ;
        RECT 58.852 61.39 75.78 61.478 ;
        RECT 59.864 60.378 76.817 60.441 ;
        RECT 75.734 44.508 75.78 61.478 ;
        RECT 58.806 61.436 75.734 61.524 ;
        RECT 59.91 60.332 76.863 60.395 ;
        RECT 75.688 44.554 75.734 61.524 ;
        RECT 58.76 61.482 75.688 61.57 ;
        RECT 59.956 60.286 76.909 60.349 ;
      LAYER MET2 ;
        RECT 70.814 69.423 79.278 69.485 ;
        RECT 77.852 62.385 110 63.5 ;
        RECT 79.232 61.005 79.278 69.485 ;
        RECT 70.768 69.469 79.232 69.531 ;
        RECT 77.898 62.339 110 63.5 ;
        RECT 79.186 61.051 79.232 69.531 ;
        RECT 70.722 69.515 79.186 69.577 ;
        RECT 77.944 62.293 110 63.5 ;
        RECT 79.14 61.097 79.186 69.577 ;
        RECT 70.676 69.561 79.14 69.623 ;
        RECT 77.99 62.247 110 63.5 ;
        RECT 79.094 61.143 79.14 69.623 ;
        RECT 70.63 69.607 79.094 69.669 ;
        RECT 78.036 62.201 110 63.5 ;
        RECT 79.048 61.189 79.094 69.669 ;
        RECT 70.584 69.653 79.048 69.715 ;
        RECT 78.082 62.155 110 63.5 ;
        RECT 79.002 61.235 79.048 69.715 ;
        RECT 70.538 69.699 79.002 69.761 ;
        RECT 78.128 62.109 110 63.5 ;
        RECT 78.956 61.281 79.002 69.761 ;
        RECT 70.492 69.745 78.956 69.807 ;
        RECT 78.174 62.063 110 63.5 ;
        RECT 78.91 61.327 78.956 69.807 ;
        RECT 70.446 69.791 78.91 69.853 ;
        RECT 78.22 62.017 110 63.5 ;
        RECT 78.864 61.373 78.91 69.853 ;
        RECT 70.4 69.837 78.864 69.899 ;
        RECT 78.266 61.971 110 63.5 ;
        RECT 78.818 61.419 78.864 69.899 ;
        RECT 70.354 69.883 78.818 69.945 ;
        RECT 78.312 61.925 110 63.5 ;
        RECT 78.772 61.465 78.818 69.945 ;
        RECT 70.308 69.929 78.772 69.991 ;
        RECT 78.358 61.879 110 63.5 ;
        RECT 78.726 61.511 78.772 69.991 ;
        RECT 70.262 69.975 78.726 70.037 ;
        RECT 78.404 61.833 110 63.5 ;
        RECT 78.68 61.557 78.726 70.037 ;
        RECT 70.216 70.021 78.68 70.083 ;
        RECT 78.45 61.787 110 63.5 ;
        RECT 78.634 61.603 78.68 70.083 ;
        RECT 70.17 70.067 78.634 70.129 ;
        RECT 78.496 61.741 110 63.5 ;
        RECT 78.588 61.649 78.634 70.129 ;
        RECT 70.124 70.113 78.588 70.175 ;
        RECT 78.542 61.695 110 63.5 ;
        RECT 70.078 70.159 78.542 70.221 ;
        RECT 70.032 70.205 78.496 70.267 ;
        RECT 69.986 70.251 78.45 70.313 ;
        RECT 69.94 70.297 78.404 70.359 ;
        RECT 69.894 70.343 78.358 70.405 ;
        RECT 69.848 70.389 78.312 70.451 ;
        RECT 69.802 70.435 78.266 70.497 ;
        RECT 69.756 70.481 78.22 70.543 ;
        RECT 69.71 70.527 78.174 70.589 ;
        RECT 69.664 70.573 78.128 70.635 ;
        RECT 69.618 70.619 78.082 70.681 ;
        RECT 69.572 70.665 78.036 70.727 ;
        RECT 69.526 70.711 77.99 70.773 ;
        RECT 69.48 70.757 77.944 70.819 ;
        RECT 69.434 70.803 77.898 70.865 ;
        RECT 69.388 70.849 77.852 70.911 ;
        RECT 69.342 70.895 77.806 70.957 ;
        RECT 69.296 70.941 77.76 71.003 ;
        RECT 69.25 70.987 77.714 71.049 ;
        RECT 69.204 71.033 77.668 71.095 ;
        RECT 69.158 71.079 77.622 71.141 ;
        RECT 69.112 71.125 77.576 71.187 ;
        RECT 69.066 71.171 77.53 71.233 ;
        RECT 69.02 71.217 77.484 71.279 ;
        RECT 68.974 71.263 77.438 71.325 ;
        RECT 68.928 71.309 77.392 71.371 ;
        RECT 68.882 71.355 77.346 71.417 ;
        RECT 68.836 71.401 77.3 71.463 ;
        RECT 68.79 71.447 77.254 71.509 ;
        RECT 68.744 71.493 77.208 71.555 ;
        RECT 68.698 71.539 77.162 71.601 ;
        RECT 68.652 71.585 77.116 71.647 ;
        RECT 68.606 71.631 77.07 71.693 ;
        RECT 68.56 71.677 77.024 71.739 ;
        RECT 68.514 71.723 76.978 71.785 ;
        RECT 68.468 71.769 76.932 71.831 ;
        RECT 68.422 71.815 76.886 71.877 ;
        RECT 68.376 71.861 76.84 71.923 ;
        RECT 68.33 71.907 76.794 71.969 ;
        RECT 68.284 71.953 76.748 72.015 ;
        RECT 68.238 71.999 76.702 72.061 ;
        RECT 68.192 72.045 76.656 72.107 ;
        RECT 68.146 72.091 76.61 72.153 ;
        RECT 68.1 72.137 76.564 72.199 ;
        RECT 68.054 72.183 76.518 72.245 ;
        RECT 68.008 72.229 76.472 72.291 ;
        RECT 67.962 72.275 76.426 72.337 ;
        RECT 67.916 72.321 76.38 72.383 ;
        RECT 67.87 72.367 76.334 72.429 ;
        RECT 67.824 72.413 76.288 72.475 ;
        RECT 67.778 72.459 76.242 72.521 ;
        RECT 67.732 72.505 76.196 72.567 ;
        RECT 67.686 72.551 76.15 72.613 ;
        RECT 67.64 72.597 76.104 72.659 ;
        RECT 67.594 72.643 76.058 72.705 ;
        RECT 67.548 72.689 76.012 72.751 ;
        RECT 67.502 72.735 75.966 72.797 ;
        RECT 67.456 72.781 75.92 72.843 ;
        RECT 67.41 72.827 75.874 72.889 ;
        RECT 67.364 72.873 75.828 72.935 ;
        RECT 67.318 72.919 75.782 72.981 ;
        RECT 67.272 72.965 75.736 73.027 ;
        RECT 67.226 73.011 75.69 73.073 ;
        RECT 67.18 73.057 75.644 73.119 ;
        RECT 67.134 73.103 75.598 73.165 ;
        RECT 67.088 73.149 75.552 73.211 ;
        RECT 67.042 73.195 75.506 73.257 ;
        RECT 66.996 73.241 75.46 73.303 ;
        RECT 66.95 73.287 75.414 73.349 ;
        RECT 66.904 73.333 75.368 73.395 ;
        RECT 66.858 73.379 75.322 73.441 ;
        RECT 66.812 73.425 75.276 73.487 ;
        RECT 66.766 73.471 75.23 73.533 ;
        RECT 66.72 73.517 75.184 73.579 ;
        RECT 66.674 73.563 75.138 73.625 ;
        RECT 66.628 73.609 75.092 73.671 ;
        RECT 66.582 73.655 75.046 73.717 ;
        RECT 66.536 73.701 75 73.763 ;
        RECT 66.49 73.747 74.954 73.809 ;
        RECT 66.444 73.793 74.908 73.855 ;
        RECT 66.398 73.839 74.862 73.901 ;
        RECT 66.352 73.885 74.816 73.947 ;
        RECT 66.306 73.931 74.77 73.993 ;
        RECT 66.26 73.977 74.724 74.039 ;
        RECT 66.214 74.023 74.678 74.085 ;
        RECT 66.168 74.069 74.632 74.131 ;
        RECT 66.122 74.115 74.586 74.177 ;
        RECT 66.076 74.161 74.54 74.223 ;
        RECT 66.03 74.207 74.494 74.269 ;
        RECT 65.984 74.253 74.448 74.315 ;
        RECT 65.938 74.299 74.402 74.361 ;
        RECT 65.892 74.345 74.356 74.407 ;
        RECT 65.846 74.391 74.31 74.453 ;
        RECT 65.8 74.437 74.264 74.499 ;
        RECT 65.754 74.483 74.218 74.545 ;
        RECT 65.708 74.529 74.172 74.591 ;
        RECT 65.662 74.575 74.126 74.637 ;
        RECT 65.616 74.621 74.08 74.683 ;
        RECT 65.57 74.667 74.034 74.729 ;
        RECT 65.524 74.713 73.988 74.775 ;
        RECT 65.478 74.759 73.942 74.821 ;
        RECT 65.432 74.805 73.896 74.867 ;
        RECT 65.386 74.851 73.85 74.913 ;
        RECT 65.34 74.897 73.804 74.959 ;
        RECT 65.294 74.943 73.758 75.005 ;
        RECT 65.248 74.989 73.712 75.051 ;
        RECT 65.202 75.035 73.666 75.097 ;
        RECT 65.156 75.081 73.62 75.143 ;
        RECT 65.11 75.127 73.574 75.189 ;
        RECT 65.064 75.173 73.528 75.235 ;
        RECT 65.018 75.219 73.482 75.281 ;
        RECT 64.972 75.265 73.436 75.327 ;
        RECT 64.926 75.311 73.39 75.373 ;
        RECT 64.88 75.357 73.344 75.419 ;
        RECT 64.834 75.403 73.298 75.465 ;
        RECT 64.788 75.449 73.252 75.511 ;
        RECT 64.742 75.495 73.206 75.557 ;
        RECT 64.696 75.541 73.16 75.603 ;
        RECT 64.65 75.587 73.114 75.649 ;
        RECT 64.604 75.633 73.068 75.695 ;
        RECT 64.558 75.679 73.022 75.741 ;
        RECT 64.512 75.725 72.976 75.787 ;
        RECT 64.466 75.771 72.93 75.833 ;
        RECT 64.42 75.817 72.884 75.879 ;
        RECT 64.374 75.863 72.838 75.925 ;
        RECT 64.328 75.909 72.792 75.971 ;
        RECT 64.282 75.955 72.746 76.017 ;
        RECT 64.236 76.001 72.7 76.063 ;
        RECT 64.19 76.047 72.654 76.109 ;
        RECT 64.144 76.093 72.608 76.155 ;
        RECT 64.098 76.139 72.562 76.201 ;
        RECT 64.052 76.185 72.516 76.247 ;
        RECT 64.006 76.231 72.47 76.293 ;
        RECT 63.96 76.277 72.424 76.339 ;
        RECT 63.914 76.323 72.378 76.385 ;
        RECT 63.868 76.369 72.332 76.431 ;
        RECT 63.822 76.415 72.286 76.477 ;
        RECT 63.776 76.461 72.24 76.523 ;
        RECT 63.73 76.507 72.194 76.569 ;
        RECT 63.684 76.553 72.148 76.615 ;
        RECT 63.638 76.599 72.102 76.661 ;
        RECT 63.592 76.645 72.056 76.707 ;
        RECT 63.546 76.691 72.01 76.753 ;
        RECT 63.5 76.737 71.964 76.799 ;
        RECT 63.48 76.77 71.918 76.845 ;
        RECT 63.434 76.803 71.872 76.891 ;
        RECT 63.388 76.849 71.826 76.937 ;
        RECT 63.342 76.895 71.78 76.983 ;
        RECT 63.296 76.941 71.734 77.029 ;
        RECT 63.25 76.987 71.688 77.075 ;
        RECT 63.204 77.033 71.642 77.121 ;
        RECT 63.158 77.079 71.596 77.167 ;
        RECT 63.112 77.125 71.55 77.213 ;
        RECT 63.066 77.171 71.504 77.259 ;
        RECT 63.02 77.217 71.458 77.305 ;
        RECT 62.974 77.263 71.412 77.351 ;
        RECT 62.928 77.309 71.366 77.397 ;
        RECT 62.882 77.355 71.32 77.443 ;
        RECT 62.836 77.401 71.274 77.489 ;
        RECT 62.79 77.447 71.228 77.535 ;
        RECT 62.744 77.493 71.182 77.581 ;
        RECT 62.698 77.539 71.136 77.627 ;
        RECT 62.652 77.585 71.09 77.673 ;
        RECT 62.606 77.631 71.044 77.719 ;
        RECT 62.56 77.677 70.998 77.765 ;
        RECT 62.514 77.723 70.952 77.811 ;
        RECT 62.468 77.769 70.906 77.857 ;
        RECT 62.422 77.815 70.86 77.903 ;
        RECT 62.376 77.861 70.814 77.949 ;
        RECT 62.33 77.907 70.768 77.995 ;
        RECT 62.284 77.953 70.722 78.041 ;
        RECT 62.238 77.999 70.676 78.087 ;
        RECT 62.192 78.045 70.63 78.133 ;
        RECT 62.146 78.091 70.584 78.179 ;
        RECT 62.1 78.137 70.538 78.225 ;
        RECT 62.054 78.183 70.492 78.271 ;
        RECT 62.008 78.229 70.446 78.317 ;
        RECT 61.962 78.275 70.4 78.363 ;
        RECT 61.916 78.321 70.354 78.409 ;
        RECT 61.87 78.367 70.308 78.455 ;
        RECT 61.824 78.413 70.262 78.501 ;
        RECT 61.778 78.459 70.216 78.547 ;
        RECT 61.732 78.505 70.17 78.593 ;
        RECT 61.686 78.551 70.124 78.639 ;
        RECT 61.64 78.597 70.078 78.685 ;
        RECT 61.594 78.643 70.032 78.731 ;
        RECT 61.548 78.689 69.986 78.777 ;
        RECT 61.502 78.735 69.94 78.823 ;
        RECT 61.456 78.781 69.894 78.869 ;
        RECT 61.41 78.827 69.848 78.915 ;
        RECT 61.364 78.873 69.802 78.961 ;
        RECT 61.318 78.919 69.756 79.007 ;
        RECT 61.272 78.965 69.71 79.053 ;
        RECT 61.226 79.011 69.664 79.099 ;
        RECT 61.18 79.057 69.618 79.145 ;
        RECT 61.134 79.103 69.572 79.191 ;
        RECT 61.088 79.149 69.526 79.237 ;
        RECT 61.042 79.195 69.48 79.283 ;
        RECT 60.996 79.241 69.434 79.329 ;
        RECT 60.95 79.287 69.388 79.375 ;
        RECT 60.904 79.333 69.342 79.421 ;
        RECT 60.858 79.379 69.296 79.467 ;
        RECT 60.812 79.425 69.25 79.513 ;
        RECT 60.766 79.471 69.204 79.559 ;
        RECT 60.72 79.517 69.158 79.605 ;
        RECT 60.674 79.563 69.112 79.651 ;
        RECT 60.628 79.609 69.066 79.697 ;
        RECT 60.582 79.655 69.02 79.743 ;
        RECT 60.536 79.701 68.974 79.789 ;
        RECT 60.49 79.747 68.928 79.835 ;
        RECT 60.444 79.793 68.882 79.881 ;
        RECT 60.398 79.839 68.836 79.927 ;
        RECT 60.352 79.885 68.79 79.973 ;
        RECT 60.306 79.931 68.744 80.019 ;
        RECT 60.26 79.977 68.698 80.065 ;
        RECT 60.214 80.023 68.652 80.111 ;
        RECT 60.168 80.069 68.606 80.157 ;
        RECT 60.122 80.115 68.56 80.203 ;
        RECT 60.076 80.161 68.514 80.249 ;
        RECT 60.03 80.207 68.468 80.295 ;
        RECT 59.984 80.253 68.422 80.341 ;
        RECT 59.938 80.299 68.376 80.387 ;
        RECT 59.892 80.345 68.33 80.433 ;
        RECT 59.846 80.391 68.284 80.479 ;
        RECT 59.8 80.437 68.238 80.525 ;
        RECT 59.754 80.483 68.192 80.571 ;
        RECT 59.708 80.529 68.146 80.617 ;
        RECT 59.662 80.575 68.1 80.663 ;
        RECT 59.616 80.621 68.054 80.709 ;
        RECT 59.57 80.667 68.008 80.755 ;
        RECT 59.524 80.713 67.962 80.801 ;
        RECT 59.478 80.759 67.916 80.847 ;
        RECT 59.432 80.805 67.87 80.893 ;
        RECT 59.386 80.851 67.824 80.939 ;
        RECT 59.34 80.897 67.778 80.985 ;
        RECT 59.294 80.943 67.732 81.031 ;
        RECT 59.248 80.989 67.686 81.077 ;
        RECT 59.202 81.035 67.64 81.123 ;
        RECT 59.156 81.081 67.594 81.169 ;
        RECT 59.11 81.127 67.548 81.215 ;
        RECT 59.064 81.173 67.502 81.261 ;
        RECT 59.018 81.219 67.456 81.307 ;
        RECT 58.972 81.265 67.41 81.353 ;
        RECT 58.926 81.311 67.364 81.399 ;
        RECT 58.88 81.357 67.318 81.445 ;
        RECT 58.834 81.403 67.272 81.491 ;
        RECT 58.788 81.449 67.226 81.537 ;
        RECT 58.742 81.495 67.18 81.583 ;
        RECT 58.696 81.541 67.134 81.629 ;
        RECT 58.65 81.587 67.088 81.675 ;
        RECT 58.604 81.633 67.042 81.721 ;
        RECT 58.558 81.679 66.996 81.767 ;
        RECT 58.512 81.725 66.95 81.813 ;
        RECT 58.466 81.771 66.904 81.859 ;
        RECT 58.42 81.817 66.858 81.905 ;
        RECT 58.374 81.863 66.812 81.951 ;
        RECT 58.328 81.909 66.766 81.997 ;
        RECT 58.282 81.955 66.72 82.043 ;
        RECT 58.236 82.001 66.674 82.089 ;
        RECT 58.19 82.047 66.628 82.135 ;
        RECT 58.144 82.093 66.582 82.181 ;
        RECT 58.098 82.139 66.536 82.227 ;
        RECT 58.052 82.185 66.49 82.273 ;
        RECT 58.006 82.231 66.444 82.319 ;
        RECT 57.96 82.277 66.398 82.365 ;
        RECT 57.914 82.323 66.352 82.411 ;
        RECT 57.868 82.369 66.306 82.457 ;
        RECT 57.822 82.415 66.26 82.503 ;
        RECT 57.776 82.461 66.214 82.549 ;
        RECT 57.73 82.507 66.168 82.595 ;
        RECT 57.684 82.553 66.122 82.641 ;
        RECT 57.638 82.599 66.076 82.687 ;
        RECT 57.592 82.645 66.03 82.733 ;
        RECT 57.546 82.691 65.984 82.779 ;
        RECT 57.5 82.737 65.938 82.825 ;
        RECT 57.5 82.737 65.892 82.871 ;
        RECT 57.5 82.737 65.846 82.917 ;
        RECT 57.5 82.737 65.8 82.963 ;
        RECT 57.5 82.737 65.754 83.009 ;
        RECT 57.5 82.737 65.708 83.055 ;
        RECT 57.5 82.737 65.662 83.101 ;
        RECT 57.5 82.737 65.616 83.147 ;
        RECT 57.5 82.737 65.57 83.193 ;
        RECT 57.5 82.737 65.524 83.239 ;
        RECT 57.5 82.737 65.478 83.285 ;
        RECT 57.5 82.737 65.432 83.331 ;
        RECT 57.5 82.737 65.386 83.377 ;
        RECT 57.5 82.737 65.34 83.423 ;
        RECT 57.5 82.737 65.294 83.469 ;
        RECT 57.5 82.737 65.248 83.515 ;
        RECT 57.5 82.737 65.202 83.561 ;
        RECT 57.5 82.737 65.156 83.607 ;
        RECT 57.5 82.737 65.11 83.653 ;
        RECT 57.5 82.737 65.064 83.699 ;
        RECT 57.5 82.737 65.018 83.745 ;
        RECT 57.5 82.737 64.972 83.791 ;
        RECT 57.5 82.737 64.926 83.837 ;
        RECT 57.5 82.737 64.88 83.883 ;
        RECT 57.5 82.737 64.834 83.929 ;
        RECT 57.5 82.737 64.788 83.975 ;
        RECT 57.5 82.737 64.742 84.021 ;
        RECT 57.5 82.737 64.696 84.067 ;
        RECT 57.5 82.737 64.65 84.113 ;
        RECT 57.5 82.737 64.604 84.159 ;
        RECT 57.5 82.737 64.558 84.205 ;
        RECT 57.5 82.737 64.512 84.251 ;
        RECT 57.5 82.737 64.466 84.297 ;
        RECT 57.5 82.737 64.42 84.343 ;
        RECT 57.5 82.737 64.374 84.389 ;
        RECT 57.5 82.737 64.328 84.435 ;
        RECT 57.5 82.737 64.282 84.481 ;
        RECT 57.5 82.737 64.236 84.527 ;
        RECT 57.5 82.737 64.19 84.573 ;
        RECT 57.5 82.737 64.144 84.619 ;
        RECT 57.5 82.737 64.098 84.665 ;
        RECT 57.5 82.737 64.052 84.711 ;
        RECT 57.5 82.737 64.006 84.757 ;
        RECT 57.5 82.737 63.96 84.803 ;
        RECT 57.5 82.737 63.914 84.849 ;
        RECT 57.5 82.737 63.868 84.895 ;
        RECT 57.5 82.737 63.822 84.941 ;
        RECT 57.5 82.737 63.776 84.987 ;
        RECT 57.5 82.737 63.73 85.033 ;
        RECT 57.5 82.737 63.684 85.079 ;
        RECT 57.5 82.737 63.638 85.125 ;
        RECT 57.5 82.737 63.592 85.171 ;
        RECT 57.5 82.737 63.546 85.217 ;
        RECT 57.5 82.737 63.5 110 ;
        RECT 88.365 68.5 110 77 ;
        RECT 79.852 76.99 91.885 77.012 ;
        RECT 76.366 80.476 88.365 80.522 ;
        RECT 76.412 80.43 88.411 80.497 ;
        RECT 88.362 68.501 88.365 80.522 ;
        RECT 76.458 80.384 88.457 80.451 ;
        RECT 88.316 68.526 88.362 80.546 ;
        RECT 76.32 80.522 88.316 80.592 ;
        RECT 76.504 80.338 88.503 80.405 ;
        RECT 88.27 68.572 88.316 80.592 ;
        RECT 76.274 80.568 88.27 80.638 ;
        RECT 76.55 80.292 88.549 80.359 ;
        RECT 88.224 68.618 88.27 80.638 ;
        RECT 76.228 80.614 88.224 80.684 ;
        RECT 76.596 80.246 88.595 80.313 ;
        RECT 88.178 68.664 88.224 80.684 ;
        RECT 76.182 80.66 88.178 80.73 ;
        RECT 76.642 80.2 88.641 80.267 ;
        RECT 88.132 68.71 88.178 80.73 ;
        RECT 76.136 80.706 88.132 80.776 ;
        RECT 76.688 80.154 88.687 80.221 ;
        RECT 88.086 68.756 88.132 80.776 ;
        RECT 76.09 80.752 88.086 80.822 ;
        RECT 76.734 80.108 88.733 80.175 ;
        RECT 88.04 68.802 88.086 80.822 ;
        RECT 76.044 80.798 88.04 80.868 ;
        RECT 76.78 80.062 88.779 80.129 ;
        RECT 87.994 68.848 88.04 80.868 ;
        RECT 75.998 80.844 87.994 80.914 ;
        RECT 76.826 80.016 88.825 80.083 ;
        RECT 87.948 68.894 87.994 80.914 ;
        RECT 75.952 80.89 87.948 80.96 ;
        RECT 76.872 79.97 88.871 80.037 ;
        RECT 87.902 68.94 87.948 80.96 ;
        RECT 75.906 80.936 87.902 81.006 ;
        RECT 76.918 79.924 88.917 79.991 ;
        RECT 87.856 68.986 87.902 81.006 ;
        RECT 75.86 80.982 87.856 81.052 ;
        RECT 76.964 79.883 88.963 79.945 ;
        RECT 87.81 69.032 87.856 81.052 ;
        RECT 75.814 81.028 87.81 81.098 ;
        RECT 77 79.842 89.009 79.899 ;
        RECT 87.764 69.078 87.81 81.098 ;
        RECT 75.768 81.074 87.764 81.144 ;
        RECT 77.046 79.796 89.055 79.853 ;
        RECT 87.718 69.124 87.764 81.144 ;
        RECT 75.722 81.12 87.718 81.19 ;
        RECT 77.092 79.75 89.101 79.807 ;
        RECT 87.672 69.17 87.718 81.19 ;
        RECT 75.676 81.166 87.672 81.236 ;
        RECT 77.138 79.704 89.147 79.761 ;
        RECT 87.626 69.216 87.672 81.236 ;
        RECT 75.63 81.212 87.626 81.282 ;
        RECT 77.184 79.658 89.193 79.715 ;
        RECT 87.58 69.262 87.626 81.282 ;
        RECT 75.584 81.258 87.58 81.328 ;
        RECT 77.23 79.612 89.239 79.669 ;
        RECT 87.534 69.308 87.58 81.328 ;
        RECT 75.538 81.304 87.534 81.374 ;
        RECT 77.276 79.566 89.285 79.623 ;
        RECT 87.488 69.354 87.534 81.374 ;
        RECT 75.492 81.35 87.488 81.42 ;
        RECT 77.322 79.52 89.331 79.577 ;
        RECT 87.442 69.4 87.488 81.42 ;
        RECT 75.446 81.396 87.442 81.466 ;
        RECT 77.368 79.474 89.377 79.531 ;
        RECT 87.396 69.446 87.442 81.466 ;
        RECT 75.4 81.442 87.396 81.512 ;
        RECT 77.414 79.428 89.423 79.485 ;
        RECT 87.35 69.492 87.396 81.512 ;
        RECT 75.354 81.488 87.35 81.558 ;
        RECT 77.46 79.382 89.469 79.439 ;
        RECT 87.304 69.538 87.35 81.558 ;
        RECT 75.308 81.534 87.304 81.604 ;
        RECT 77.506 79.336 89.515 79.393 ;
        RECT 87.258 69.584 87.304 81.604 ;
        RECT 75.262 81.58 87.258 81.65 ;
        RECT 77.552 79.29 89.561 79.347 ;
        RECT 87.212 69.63 87.258 81.65 ;
        RECT 75.216 81.626 87.212 81.696 ;
        RECT 77.598 79.244 89.607 79.301 ;
        RECT 87.166 69.676 87.212 81.696 ;
        RECT 75.17 81.672 87.166 81.742 ;
        RECT 77.644 79.198 89.653 79.255 ;
        RECT 87.12 69.722 87.166 81.742 ;
        RECT 75.124 81.718 87.12 81.788 ;
        RECT 77.69 79.152 89.699 79.209 ;
        RECT 87.074 69.768 87.12 81.788 ;
        RECT 75.078 81.764 87.074 81.834 ;
        RECT 77.736 79.106 89.745 79.163 ;
        RECT 87.028 69.814 87.074 81.834 ;
        RECT 75.032 81.81 87.028 81.88 ;
        RECT 77.782 79.06 89.791 79.117 ;
        RECT 86.982 69.86 87.028 81.88 ;
        RECT 74.986 81.856 86.982 81.926 ;
        RECT 77.828 79.014 89.837 79.071 ;
        RECT 86.936 69.906 86.982 81.926 ;
        RECT 74.94 81.902 86.936 81.972 ;
        RECT 77.874 78.968 89.883 79.025 ;
        RECT 86.89 69.952 86.936 81.972 ;
        RECT 74.894 81.948 86.89 82.018 ;
        RECT 77.92 78.922 89.929 78.979 ;
        RECT 86.844 69.998 86.89 82.018 ;
        RECT 74.848 81.994 86.844 82.064 ;
        RECT 77.966 78.876 89.975 78.933 ;
        RECT 86.798 70.044 86.844 82.064 ;
        RECT 74.802 82.04 86.798 82.11 ;
        RECT 78.012 78.83 90.021 78.887 ;
        RECT 86.752 70.09 86.798 82.11 ;
        RECT 74.756 82.086 86.752 82.156 ;
        RECT 78.058 78.784 90.067 78.841 ;
        RECT 86.706 70.136 86.752 82.156 ;
        RECT 74.71 82.132 86.706 82.202 ;
        RECT 78.104 78.738 90.113 78.795 ;
        RECT 86.66 70.182 86.706 82.202 ;
        RECT 74.664 82.178 86.66 82.248 ;
        RECT 78.15 78.692 90.159 78.749 ;
        RECT 86.614 70.228 86.66 82.248 ;
        RECT 74.618 82.224 86.614 82.294 ;
        RECT 78.196 78.646 90.205 78.703 ;
        RECT 86.568 70.274 86.614 82.294 ;
        RECT 74.572 82.27 86.568 82.34 ;
        RECT 78.242 78.6 90.251 78.657 ;
        RECT 86.522 70.32 86.568 82.34 ;
        RECT 74.526 82.316 86.522 82.386 ;
        RECT 78.288 78.554 90.297 78.611 ;
        RECT 86.476 70.366 86.522 82.386 ;
        RECT 74.48 82.362 86.476 82.432 ;
        RECT 78.334 78.508 90.343 78.565 ;
        RECT 86.43 70.412 86.476 82.432 ;
        RECT 74.434 82.408 86.43 82.478 ;
        RECT 78.38 78.462 90.389 78.519 ;
        RECT 86.384 70.458 86.43 82.478 ;
        RECT 74.388 82.454 86.384 82.524 ;
        RECT 78.426 78.416 90.435 78.473 ;
        RECT 86.338 70.504 86.384 82.524 ;
        RECT 74.342 82.5 86.338 82.57 ;
        RECT 78.472 78.37 90.481 78.427 ;
        RECT 86.292 70.55 86.338 82.57 ;
        RECT 74.296 82.546 86.292 82.616 ;
        RECT 78.518 78.324 90.527 78.381 ;
        RECT 86.246 70.596 86.292 82.616 ;
        RECT 74.25 82.592 86.246 82.662 ;
        RECT 78.564 78.278 90.573 78.335 ;
        RECT 86.2 70.642 86.246 82.662 ;
        RECT 74.204 82.638 86.2 82.708 ;
        RECT 78.61 78.232 90.619 78.289 ;
        RECT 86.154 70.688 86.2 82.708 ;
        RECT 74.158 82.684 86.154 82.754 ;
        RECT 78.656 78.186 90.665 78.243 ;
        RECT 86.108 70.734 86.154 82.754 ;
        RECT 74.112 82.73 86.108 82.8 ;
        RECT 78.702 78.14 90.711 78.197 ;
        RECT 86.062 70.78 86.108 82.8 ;
        RECT 74.066 82.776 86.062 82.846 ;
        RECT 78.748 78.094 90.757 78.151 ;
        RECT 86.016 70.826 86.062 82.846 ;
        RECT 74.02 82.822 86.016 82.892 ;
        RECT 78.794 78.048 90.803 78.105 ;
        RECT 85.97 70.872 86.016 82.892 ;
        RECT 73.974 82.868 85.97 82.938 ;
        RECT 78.84 78.002 90.849 78.059 ;
        RECT 85.924 70.918 85.97 82.938 ;
        RECT 73.928 82.914 85.924 82.984 ;
        RECT 78.886 77.956 90.895 78.013 ;
        RECT 85.878 70.964 85.924 82.984 ;
        RECT 73.882 82.96 85.878 83.03 ;
        RECT 78.932 77.91 90.941 77.967 ;
        RECT 85.832 71.01 85.878 83.03 ;
        RECT 73.836 83.006 85.832 83.076 ;
        RECT 78.978 77.864 90.987 77.921 ;
        RECT 85.786 71.056 85.832 83.076 ;
        RECT 73.79 83.052 85.786 83.122 ;
        RECT 79.024 77.818 91.033 77.875 ;
        RECT 85.74 71.102 85.786 83.122 ;
        RECT 73.744 83.098 85.74 83.168 ;
        RECT 79.07 77.772 91.079 77.829 ;
        RECT 85.694 71.148 85.74 83.168 ;
        RECT 73.698 83.144 85.694 83.214 ;
        RECT 79.116 77.726 91.125 77.783 ;
        RECT 85.648 71.194 85.694 83.214 ;
        RECT 73.652 83.19 85.648 83.26 ;
        RECT 79.162 77.68 91.171 77.737 ;
        RECT 85.602 71.24 85.648 83.26 ;
        RECT 73.606 83.236 85.602 83.306 ;
        RECT 79.208 77.634 91.217 77.691 ;
        RECT 85.556 71.286 85.602 83.306 ;
        RECT 73.56 83.282 85.556 83.352 ;
        RECT 79.254 77.588 91.263 77.645 ;
        RECT 85.51 71.332 85.556 83.352 ;
        RECT 73.514 83.328 85.51 83.398 ;
        RECT 79.3 77.542 91.309 77.599 ;
        RECT 85.464 71.378 85.51 83.398 ;
        RECT 73.468 83.374 85.464 83.444 ;
        RECT 79.346 77.496 91.355 77.553 ;
        RECT 85.418 71.424 85.464 83.444 ;
        RECT 73.422 83.42 85.418 83.49 ;
        RECT 79.392 77.45 91.401 77.507 ;
        RECT 85.372 71.47 85.418 83.49 ;
        RECT 73.376 83.466 85.372 83.536 ;
        RECT 79.438 77.404 91.447 77.461 ;
        RECT 85.326 71.516 85.372 83.536 ;
        RECT 73.33 83.512 85.326 83.582 ;
        RECT 79.484 77.358 91.493 77.415 ;
        RECT 85.28 71.562 85.326 83.582 ;
        RECT 73.284 83.558 85.28 83.628 ;
        RECT 79.53 77.312 91.539 77.369 ;
        RECT 85.234 71.608 85.28 83.628 ;
        RECT 73.238 83.604 85.234 83.674 ;
        RECT 79.576 77.266 91.585 77.323 ;
        RECT 85.188 71.654 85.234 83.674 ;
        RECT 73.192 83.65 85.188 83.72 ;
        RECT 79.622 77.22 91.631 77.277 ;
        RECT 85.142 71.7 85.188 83.72 ;
        RECT 73.146 83.696 85.142 83.766 ;
        RECT 79.668 77.174 91.677 77.231 ;
        RECT 85.096 71.746 85.142 83.766 ;
        RECT 73.1 83.742 85.096 83.812 ;
        RECT 79.714 77.128 91.723 77.185 ;
        RECT 85.05 71.792 85.096 83.812 ;
        RECT 73.054 83.788 85.05 83.858 ;
        RECT 79.76 77.082 91.769 77.139 ;
        RECT 85.004 71.838 85.05 83.858 ;
        RECT 73.008 83.834 85.004 83.904 ;
        RECT 79.806 77.036 91.815 77.093 ;
        RECT 84.958 71.884 85.004 83.904 ;
        RECT 72.962 83.88 84.958 83.95 ;
        RECT 79.852 76.99 91.861 77.047 ;
        RECT 84.912 71.93 84.958 83.95 ;
        RECT 72.916 83.926 84.912 83.996 ;
        RECT 79.898 76.944 110 77 ;
        RECT 84.866 71.976 84.912 83.996 ;
        RECT 72.87 83.972 84.866 84.042 ;
        RECT 79.944 76.898 110 77 ;
        RECT 84.82 72.022 84.866 84.042 ;
        RECT 72.824 84.018 84.82 84.088 ;
        RECT 79.99 76.852 110 77 ;
        RECT 84.774 72.068 84.82 84.088 ;
        RECT 72.778 84.064 84.774 84.134 ;
        RECT 80.036 76.806 110 77 ;
        RECT 84.728 72.114 84.774 84.134 ;
        RECT 72.732 84.11 84.728 84.18 ;
        RECT 80.082 76.76 110 77 ;
        RECT 84.682 72.16 84.728 84.18 ;
        RECT 72.686 84.156 84.682 84.226 ;
        RECT 80.128 76.714 110 77 ;
        RECT 84.636 72.206 84.682 84.226 ;
        RECT 72.64 84.202 84.636 84.272 ;
        RECT 80.174 76.668 110 77 ;
        RECT 84.59 72.252 84.636 84.272 ;
        RECT 72.594 84.248 84.59 84.318 ;
        RECT 80.22 76.622 110 77 ;
        RECT 84.544 72.298 84.59 84.318 ;
        RECT 72.548 84.294 84.544 84.364 ;
        RECT 80.266 76.576 110 77 ;
        RECT 84.498 72.344 84.544 84.364 ;
        RECT 72.502 84.34 84.498 84.41 ;
        RECT 80.312 76.53 110 77 ;
        RECT 84.452 72.39 84.498 84.41 ;
        RECT 72.456 84.386 84.452 84.456 ;
        RECT 80.358 76.484 110 77 ;
        RECT 84.406 72.436 84.452 84.456 ;
        RECT 72.41 84.432 84.406 84.502 ;
        RECT 80.404 76.438 110 77 ;
        RECT 84.36 72.482 84.406 84.502 ;
        RECT 72.364 84.478 84.36 84.548 ;
        RECT 80.45 76.392 110 77 ;
        RECT 84.314 72.528 84.36 84.548 ;
        RECT 72.318 84.524 84.314 84.594 ;
        RECT 80.496 76.346 110 77 ;
        RECT 84.268 72.574 84.314 84.594 ;
        RECT 72.272 84.57 84.268 84.64 ;
        RECT 80.542 76.3 110 77 ;
        RECT 84.222 72.62 84.268 84.64 ;
        RECT 72.226 84.616 84.222 84.686 ;
        RECT 80.588 76.254 110 77 ;
        RECT 84.176 72.666 84.222 84.686 ;
        RECT 72.18 84.662 84.176 84.732 ;
        RECT 80.634 76.208 110 77 ;
        RECT 84.13 72.712 84.176 84.732 ;
        RECT 72.134 84.708 84.13 84.778 ;
        RECT 80.68 76.162 110 77 ;
        RECT 84.084 72.758 84.13 84.778 ;
        RECT 72.088 84.754 84.084 84.824 ;
        RECT 80.726 76.116 110 77 ;
        RECT 84.038 72.804 84.084 84.824 ;
        RECT 72.042 84.8 84.038 84.87 ;
        RECT 80.772 76.07 110 77 ;
        RECT 83.992 72.85 84.038 84.87 ;
        RECT 71.996 84.846 83.992 84.916 ;
        RECT 80.818 76.024 110 77 ;
        RECT 83.946 72.896 83.992 84.916 ;
        RECT 71.95 84.892 83.946 84.962 ;
        RECT 80.864 75.978 110 77 ;
        RECT 83.9 72.942 83.946 84.962 ;
        RECT 71.904 84.938 83.9 85.008 ;
        RECT 80.91 75.932 110 77 ;
        RECT 83.854 72.988 83.9 85.008 ;
        RECT 71.858 84.984 83.854 85.054 ;
        RECT 80.956 75.886 110 77 ;
        RECT 83.808 73.034 83.854 85.054 ;
        RECT 71.812 85.03 83.808 85.1 ;
        RECT 81.002 75.84 110 77 ;
        RECT 83.762 73.08 83.808 85.1 ;
        RECT 71.766 85.076 83.762 85.146 ;
        RECT 81.048 75.794 110 77 ;
        RECT 83.716 73.126 83.762 85.146 ;
        RECT 71.72 85.122 83.716 85.192 ;
        RECT 81.094 75.748 110 77 ;
        RECT 83.67 73.172 83.716 85.192 ;
        RECT 71.674 85.168 83.67 85.238 ;
        RECT 81.14 75.702 110 77 ;
        RECT 83.624 73.218 83.67 85.238 ;
        RECT 71.628 85.214 83.624 85.284 ;
        RECT 81.186 75.656 110 77 ;
        RECT 83.578 73.264 83.624 85.284 ;
        RECT 71.582 85.26 83.578 85.33 ;
        RECT 81.232 75.61 110 77 ;
        RECT 83.532 73.31 83.578 85.33 ;
        RECT 71.536 85.306 83.532 85.376 ;
        RECT 81.278 75.564 110 77 ;
        RECT 83.486 73.356 83.532 85.376 ;
        RECT 71.49 85.352 83.486 85.422 ;
        RECT 81.324 75.518 110 77 ;
        RECT 83.44 73.402 83.486 85.422 ;
        RECT 71.444 85.398 83.44 85.468 ;
        RECT 81.37 75.472 110 77 ;
        RECT 83.394 73.448 83.44 85.468 ;
        RECT 71.398 85.444 83.394 85.514 ;
        RECT 81.416 75.426 110 77 ;
        RECT 83.348 73.494 83.394 85.514 ;
        RECT 71.352 85.49 83.348 85.56 ;
        RECT 81.462 75.38 110 77 ;
        RECT 83.302 73.54 83.348 85.56 ;
        RECT 71.306 85.536 83.302 85.606 ;
        RECT 81.508 75.334 110 77 ;
        RECT 83.256 73.586 83.302 85.606 ;
        RECT 71.26 85.582 83.256 85.652 ;
        RECT 81.554 75.288 110 77 ;
        RECT 83.21 73.632 83.256 85.652 ;
        RECT 71.214 85.628 83.21 85.698 ;
        RECT 81.6 75.242 110 77 ;
        RECT 83.164 73.678 83.21 85.698 ;
        RECT 71.168 85.674 83.164 85.744 ;
        RECT 81.646 75.196 110 77 ;
        RECT 83.118 73.724 83.164 85.744 ;
        RECT 71.122 85.72 83.118 85.79 ;
        RECT 81.692 75.15 110 77 ;
        RECT 83.072 73.77 83.118 85.79 ;
        RECT 71.076 85.766 83.072 85.836 ;
        RECT 81.738 75.104 110 77 ;
        RECT 83.026 73.816 83.072 85.836 ;
        RECT 71.03 85.812 83.026 85.882 ;
        RECT 81.784 75.058 110 77 ;
        RECT 82.98 73.862 83.026 85.882 ;
        RECT 70.984 85.858 82.98 85.928 ;
        RECT 81.83 75.012 110 77 ;
        RECT 82.934 73.908 82.98 85.928 ;
        RECT 70.938 85.904 82.934 85.974 ;
        RECT 81.876 74.966 110 77 ;
        RECT 82.888 73.954 82.934 85.974 ;
        RECT 70.892 85.95 82.888 86.02 ;
        RECT 81.922 74.92 110 77 ;
        RECT 82.842 74 82.888 86.02 ;
        RECT 70.846 85.996 82.842 86.066 ;
        RECT 81.968 74.874 110 77 ;
        RECT 82.796 74.046 82.842 86.066 ;
        RECT 70.8 86.042 82.796 86.112 ;
        RECT 82.014 74.828 110 77 ;
        RECT 82.75 74.092 82.796 86.112 ;
        RECT 70.754 86.088 82.75 86.158 ;
        RECT 82.06 74.782 110 77 ;
        RECT 82.704 74.138 82.75 86.158 ;
        RECT 70.708 86.134 82.704 86.204 ;
        RECT 82.106 74.736 110 77 ;
        RECT 82.658 74.184 82.704 86.204 ;
        RECT 70.662 86.18 82.658 86.25 ;
        RECT 82.152 74.69 110 77 ;
        RECT 82.612 74.23 82.658 86.25 ;
        RECT 70.616 86.226 82.612 86.296 ;
        RECT 82.198 74.644 110 77 ;
        RECT 82.566 74.276 82.612 86.296 ;
        RECT 70.57 86.272 82.566 86.342 ;
        RECT 82.244 74.598 110 77 ;
        RECT 82.52 74.322 82.566 86.342 ;
        RECT 70.524 86.318 82.52 86.388 ;
        RECT 82.29 74.552 110 77 ;
        RECT 82.474 74.368 82.52 86.388 ;
        RECT 70.478 86.364 82.474 86.434 ;
        RECT 82.336 74.506 110 77 ;
        RECT 82.428 74.414 82.474 86.434 ;
        RECT 70.432 86.41 82.428 86.48 ;
        RECT 82.382 74.46 110 77 ;
        RECT 70.386 86.456 82.382 86.526 ;
        RECT 70.34 86.502 82.336 86.572 ;
        RECT 70.294 86.548 82.29 86.618 ;
        RECT 70.248 86.594 82.244 86.664 ;
        RECT 70.202 86.64 82.198 86.71 ;
        RECT 70.156 86.686 82.152 86.756 ;
        RECT 70.11 86.732 82.106 86.802 ;
        RECT 70.064 86.778 82.06 86.848 ;
        RECT 70.018 86.824 82.014 86.894 ;
        RECT 69.972 86.87 81.968 86.94 ;
        RECT 69.926 86.916 81.922 86.986 ;
        RECT 69.88 86.962 81.876 87.032 ;
        RECT 69.834 87.008 81.83 87.078 ;
        RECT 69.788 87.054 81.784 87.124 ;
        RECT 69.742 87.1 81.738 87.17 ;
        RECT 69.696 87.146 81.692 87.216 ;
        RECT 69.65 87.192 81.646 87.262 ;
        RECT 69.604 87.238 81.6 87.308 ;
        RECT 69.558 87.284 81.554 87.354 ;
        RECT 69.512 87.33 81.508 87.4 ;
        RECT 69.466 87.376 81.462 87.446 ;
        RECT 69.42 87.422 81.416 87.492 ;
        RECT 69.374 87.468 81.37 87.538 ;
        RECT 69.328 87.514 81.324 87.584 ;
        RECT 69.282 87.56 81.278 87.63 ;
        RECT 69.236 87.606 81.232 87.676 ;
        RECT 69.19 87.652 81.186 87.722 ;
        RECT 69.144 87.698 81.14 87.768 ;
        RECT 69.098 87.744 81.094 87.814 ;
        RECT 69.052 87.79 81.048 87.86 ;
        RECT 69.006 87.836 81.002 87.906 ;
        RECT 68.96 87.882 80.956 87.952 ;
        RECT 68.914 87.928 80.91 87.998 ;
        RECT 68.868 87.974 80.864 88.044 ;
        RECT 68.822 88.02 80.818 88.09 ;
        RECT 68.776 88.066 80.772 88.136 ;
        RECT 68.73 88.112 80.726 88.182 ;
        RECT 68.684 88.158 80.68 88.228 ;
        RECT 68.638 88.204 80.634 88.274 ;
        RECT 68.592 88.25 80.588 88.32 ;
        RECT 68.546 88.296 80.542 88.366 ;
        RECT 68.5 88.342 80.496 88.412 ;
        RECT 68.5 88.342 80.45 88.458 ;
        RECT 68.5 88.342 80.404 88.504 ;
        RECT 68.5 88.342 80.358 88.55 ;
        RECT 68.5 88.342 80.312 88.596 ;
        RECT 68.5 88.342 80.266 88.642 ;
        RECT 68.5 88.342 80.22 88.688 ;
        RECT 68.5 88.342 80.174 88.734 ;
        RECT 68.5 88.342 80.128 88.78 ;
        RECT 68.5 88.342 80.082 88.826 ;
        RECT 68.5 88.342 80.036 88.872 ;
        RECT 68.5 88.342 79.99 88.918 ;
        RECT 68.5 88.342 79.944 88.964 ;
        RECT 68.5 88.342 79.898 89.01 ;
        RECT 68.5 88.342 79.852 89.056 ;
        RECT 68.5 88.342 79.806 89.102 ;
        RECT 68.5 88.342 79.76 89.148 ;
        RECT 68.5 88.342 79.714 89.194 ;
        RECT 68.5 88.342 79.668 89.24 ;
        RECT 68.5 88.342 79.622 89.286 ;
        RECT 68.5 88.342 79.576 89.332 ;
        RECT 68.5 88.342 79.53 89.378 ;
        RECT 68.5 88.342 79.484 89.424 ;
        RECT 68.5 88.342 79.438 89.47 ;
        RECT 68.5 88.342 79.392 89.516 ;
        RECT 68.5 88.342 79.346 89.562 ;
        RECT 68.5 88.342 79.3 89.608 ;
        RECT 68.5 88.342 79.254 89.654 ;
        RECT 68.5 88.342 79.208 89.7 ;
        RECT 68.5 88.342 79.162 89.746 ;
        RECT 68.5 88.342 79.116 89.792 ;
        RECT 68.5 88.342 79.07 89.838 ;
        RECT 68.5 88.342 79.024 89.884 ;
        RECT 68.5 88.342 78.978 89.93 ;
        RECT 68.5 88.342 78.932 89.976 ;
        RECT 68.5 88.342 78.886 90.022 ;
        RECT 68.5 88.342 78.84 90.068 ;
        RECT 68.5 88.342 78.794 90.114 ;
        RECT 68.5 88.342 78.748 90.16 ;
        RECT 68.5 88.342 78.702 90.206 ;
        RECT 68.5 88.342 78.656 90.252 ;
        RECT 68.5 88.342 78.61 90.298 ;
        RECT 68.5 88.342 78.564 90.344 ;
        RECT 68.5 88.342 78.518 90.39 ;
        RECT 68.5 88.342 78.472 90.436 ;
        RECT 68.5 88.342 78.426 90.482 ;
        RECT 68.5 88.342 78.38 90.528 ;
        RECT 68.5 88.342 78.334 90.574 ;
        RECT 68.5 88.342 78.288 90.62 ;
        RECT 68.5 88.342 78.242 90.666 ;
        RECT 68.5 88.342 78.196 90.712 ;
        RECT 68.5 88.342 78.15 90.758 ;
        RECT 68.5 88.342 78.104 90.804 ;
        RECT 68.5 88.342 78.058 90.85 ;
        RECT 68.5 88.342 78.012 90.896 ;
        RECT 68.5 88.342 77.966 90.942 ;
        RECT 68.5 88.342 77.92 90.988 ;
        RECT 68.5 88.342 77.874 91.034 ;
        RECT 68.5 88.342 77.828 91.08 ;
        RECT 68.5 88.342 77.782 91.126 ;
        RECT 68.5 88.342 77.736 91.172 ;
        RECT 68.5 88.342 77.69 91.218 ;
        RECT 68.5 88.342 77.644 91.264 ;
        RECT 68.5 88.342 77.598 91.31 ;
        RECT 68.5 88.342 77.552 91.356 ;
        RECT 68.5 88.342 77.506 91.402 ;
        RECT 68.5 88.342 77.46 91.448 ;
        RECT 68.5 88.342 77.414 91.494 ;
        RECT 68.5 88.342 77.368 91.54 ;
        RECT 68.5 88.342 77.322 91.586 ;
        RECT 68.5 88.342 77.276 91.632 ;
        RECT 68.5 88.342 77.23 91.678 ;
        RECT 68.5 88.342 77.184 91.724 ;
        RECT 68.5 88.342 77.138 91.77 ;
        RECT 68.5 88.342 77.092 91.816 ;
        RECT 68.5 88.342 77.046 91.862 ;
        RECT 68.5 88.342 77 110 ;
        RECT 75.642 44.6 75.688 61.57 ;
        RECT 58.714 61.528 75.642 61.616 ;
        RECT 60.002 60.24 76.955 60.303 ;
        RECT 75.596 44.646 75.642 61.616 ;
        RECT 58.668 61.574 75.596 61.662 ;
        RECT 60.048 60.194 77.001 60.257 ;
        RECT 75.55 44.692 75.596 61.662 ;
        RECT 58.622 61.62 75.55 61.708 ;
        RECT 60.094 60.148 77.047 60.211 ;
        RECT 75.504 44.738 75.55 61.708 ;
        RECT 58.576 61.666 75.504 61.754 ;
        RECT 60.14 60.102 77.093 60.165 ;
        RECT 75.458 44.784 75.504 61.754 ;
        RECT 58.53 61.712 75.458 61.8 ;
        RECT 60.186 60.056 77.139 60.119 ;
        RECT 75.412 44.83 75.458 61.8 ;
        RECT 58.484 61.758 75.412 61.846 ;
        RECT 60.232 60.01 77.185 60.073 ;
        RECT 75.366 44.876 75.412 61.846 ;
        RECT 58.438 61.804 75.366 61.892 ;
        RECT 60.278 59.964 77.231 60.027 ;
        RECT 75.32 44.922 75.366 61.892 ;
        RECT 58.392 61.85 75.32 61.938 ;
        RECT 60.324 59.918 77.277 59.981 ;
        RECT 75.274 44.968 75.32 61.938 ;
        RECT 58.346 61.896 75.274 61.984 ;
        RECT 60.37 59.872 77.323 59.935 ;
        RECT 75.228 45.014 75.274 61.984 ;
        RECT 58.3 61.942 75.228 62.03 ;
        RECT 60.416 59.826 77.369 59.889 ;
        RECT 75.182 45.06 75.228 62.03 ;
        RECT 58.254 61.988 75.182 62.076 ;
        RECT 60.462 59.78 77.415 59.843 ;
        RECT 75.136 45.106 75.182 62.076 ;
        RECT 58.208 62.034 75.136 62.122 ;
        RECT 60.508 59.734 77.461 59.797 ;
        RECT 75.09 45.152 75.136 62.122 ;
        RECT 58.162 62.08 75.09 62.168 ;
        RECT 60.554 59.688 77.507 59.751 ;
        RECT 75.044 45.198 75.09 62.168 ;
        RECT 58.116 62.126 75.044 62.214 ;
        RECT 60.6 59.642 77.553 59.705 ;
        RECT 74.998 45.244 75.044 62.214 ;
        RECT 58.07 62.172 74.998 62.26 ;
        RECT 60.646 59.596 77.599 59.659 ;
        RECT 74.952 45.29 74.998 62.26 ;
        RECT 58.024 62.218 74.952 62.306 ;
        RECT 60.692 59.55 77.645 59.613 ;
        RECT 74.906 45.336 74.952 62.306 ;
        RECT 57.978 62.264 74.906 62.352 ;
        RECT 60.738 59.504 77.691 59.567 ;
        RECT 74.86 45.382 74.906 62.352 ;
        RECT 57.932 62.31 74.86 62.398 ;
        RECT 60.784 59.458 77.737 59.521 ;
        RECT 74.814 45.428 74.86 62.398 ;
        RECT 57.886 62.356 74.814 62.444 ;
        RECT 60.83 59.412 77.783 59.475 ;
        RECT 74.768 45.474 74.814 62.444 ;
        RECT 57.84 62.402 74.768 62.49 ;
        RECT 60.876 59.366 77.829 59.429 ;
        RECT 74.722 45.52 74.768 62.49 ;
        RECT 57.794 62.448 74.722 62.536 ;
        RECT 60.922 59.32 77.875 59.383 ;
        RECT 74.676 45.566 74.722 62.536 ;
        RECT 57.748 62.494 74.676 62.582 ;
        RECT 60.968 59.274 77.921 59.337 ;
        RECT 74.63 45.612 74.676 62.582 ;
        RECT 57.702 62.54 74.63 62.628 ;
        RECT 61.014 59.228 77.967 59.291 ;
        RECT 74.584 45.658 74.63 62.628 ;
        RECT 57.656 62.586 74.584 62.674 ;
        RECT 61.06 59.182 78.013 59.245 ;
        RECT 74.538 45.704 74.584 62.674 ;
        RECT 57.61 62.632 74.538 62.72 ;
        RECT 61.106 59.136 78.059 59.199 ;
        RECT 74.492 45.75 74.538 62.72 ;
        RECT 57.564 62.678 74.492 62.766 ;
        RECT 61.152 59.09 78.105 59.153 ;
        RECT 74.446 45.796 74.492 62.766 ;
        RECT 57.518 62.724 74.446 62.812 ;
        RECT 61.198 59.044 78.151 59.107 ;
        RECT 74.4 45.842 74.446 62.812 ;
        RECT 57.472 62.77 74.4 62.858 ;
        RECT 61.244 58.998 78.197 59.061 ;
        RECT 74.354 45.888 74.4 62.858 ;
        RECT 57.426 62.816 74.354 62.904 ;
        RECT 61.29 58.952 78.243 59.015 ;
        RECT 74.308 45.934 74.354 62.904 ;
        RECT 57.38 62.862 74.308 62.95 ;
        RECT 61.336 58.906 78.289 58.969 ;
        RECT 74.262 45.98 74.308 62.95 ;
        RECT 57.334 62.908 74.262 62.996 ;
        RECT 61.382 58.86 78.335 58.923 ;
        RECT 74.216 46.026 74.262 62.996 ;
        RECT 57.288 62.954 74.216 63.042 ;
        RECT 61.428 58.814 78.381 58.877 ;
        RECT 74.17 46.072 74.216 63.042 ;
        RECT 57.242 63 74.17 63.088 ;
        RECT 61.474 58.768 78.427 58.831 ;
        RECT 74.124 46.118 74.17 63.088 ;
        RECT 57.196 63.046 74.124 63.134 ;
        RECT 61.52 58.722 78.473 58.785 ;
        RECT 74.078 46.164 74.124 63.134 ;
        RECT 57.15 63.092 74.078 63.18 ;
        RECT 61.566 58.676 78.519 58.739 ;
        RECT 74.032 46.21 74.078 63.18 ;
        RECT 57.104 63.138 74.032 63.226 ;
        RECT 61.612 58.63 78.565 58.693 ;
        RECT 73.986 46.256 74.032 63.226 ;
        RECT 57.058 63.184 73.986 63.272 ;
        RECT 61.658 58.584 78.611 58.647 ;
        RECT 73.94 46.302 73.986 63.272 ;
        RECT 57.012 63.23 73.94 63.318 ;
        RECT 61.704 58.538 78.657 58.601 ;
        RECT 73.894 46.348 73.94 63.318 ;
        RECT 56.966 63.276 73.894 63.364 ;
        RECT 61.75 58.492 78.703 58.555 ;
        RECT 73.848 46.394 73.894 63.364 ;
        RECT 56.92 63.322 73.848 63.41 ;
        RECT 61.796 58.446 78.749 58.509 ;
        RECT 73.802 46.44 73.848 63.41 ;
        RECT 56.874 63.368 73.802 63.456 ;
        RECT 61.842 58.4 78.795 58.463 ;
        RECT 73.756 46.486 73.802 63.456 ;
        RECT 56.828 63.414 73.756 63.502 ;
        RECT 61.888 58.354 78.841 58.417 ;
        RECT 73.71 46.532 73.756 63.502 ;
        RECT 56.782 63.46 73.71 63.548 ;
        RECT 61.934 58.308 78.887 58.371 ;
        RECT 73.664 46.578 73.71 63.548 ;
        RECT 56.736 63.506 73.664 63.594 ;
        RECT 61.98 58.262 78.933 58.325 ;
        RECT 73.618 46.624 73.664 63.594 ;
        RECT 56.69 63.552 73.618 63.64 ;
        RECT 62.026 58.216 78.979 58.279 ;
        RECT 73.572 46.67 73.618 63.64 ;
        RECT 56.644 63.598 73.572 63.686 ;
        RECT 62.072 58.17 79.025 58.233 ;
        RECT 73.526 46.716 73.572 63.686 ;
        RECT 56.598 63.644 73.526 63.732 ;
        RECT 62.118 58.124 79.071 58.187 ;
        RECT 73.48 46.762 73.526 63.732 ;
        RECT 56.552 63.69 73.48 63.778 ;
        RECT 62.164 58.078 79.117 58.141 ;
        RECT 73.434 46.808 73.48 63.778 ;
        RECT 56.506 63.736 73.434 63.824 ;
        RECT 62.21 58.032 79.163 58.095 ;
        RECT 73.388 46.854 73.434 63.824 ;
        RECT 56.46 63.782 73.388 63.87 ;
        RECT 62.256 57.986 79.209 58.049 ;
        RECT 73.342 46.9 73.388 63.87 ;
        RECT 56.414 63.828 73.342 63.916 ;
        RECT 62.302 57.94 79.255 58.003 ;
        RECT 73.296 46.946 73.342 63.916 ;
        RECT 56.368 63.874 73.296 63.962 ;
        RECT 62.348 57.894 79.301 57.957 ;
        RECT 73.25 46.992 73.296 63.962 ;
        RECT 56.322 63.92 73.25 64.008 ;
        RECT 62.394 57.848 79.347 57.911 ;
        RECT 73.204 47.038 73.25 64.008 ;
        RECT 56.276 63.966 73.204 64.054 ;
        RECT 62.44 57.802 79.393 57.865 ;
        RECT 73.158 47.084 73.204 64.054 ;
        RECT 56.23 64.012 73.158 64.1 ;
        RECT 62.486 57.756 79.439 57.819 ;
        RECT 73.112 47.13 73.158 64.1 ;
        RECT 56.184 64.058 73.112 64.146 ;
        RECT 62.532 57.71 79.485 57.773 ;
        RECT 73.066 47.176 73.112 64.146 ;
        RECT 56.138 64.104 73.066 64.192 ;
        RECT 62.578 57.664 79.531 57.727 ;
        RECT 73.02 47.222 73.066 64.192 ;
        RECT 56.092 64.15 73.02 64.238 ;
        RECT 62.624 57.618 79.577 57.681 ;
        RECT 72.974 47.268 73.02 64.238 ;
        RECT 56 64.242 72.974 64.284 ;
        RECT 56.046 64.196 72.974 64.284 ;
        RECT 62.67 57.572 79.623 57.635 ;
        RECT 72.928 47.314 72.974 64.284 ;
        RECT 55.96 64.285 72.928 64.33 ;
        RECT 62.716 57.526 79.669 57.589 ;
        RECT 72.882 47.36 72.928 64.33 ;
        RECT 55.914 64.328 72.882 64.376 ;
        RECT 62.762 57.48 79.715 57.543 ;
        RECT 72.836 47.406 72.882 64.376 ;
        RECT 55.868 64.374 72.836 64.422 ;
        RECT 62.808 57.434 79.761 57.497 ;
        RECT 72.79 47.452 72.836 64.422 ;
        RECT 55.822 64.42 72.79 64.468 ;
        RECT 62.854 57.388 79.807 57.451 ;
        RECT 72.744 47.498 72.79 64.468 ;
        RECT 55.776 64.466 72.744 64.514 ;
        RECT 62.9 57.342 79.853 57.405 ;
        RECT 72.698 47.544 72.744 64.514 ;
        RECT 55.73 64.512 72.698 64.56 ;
        RECT 62.946 57.296 79.899 57.359 ;
        RECT 72.652 47.59 72.698 64.56 ;
        RECT 55.684 64.558 72.652 64.606 ;
        RECT 62.992 57.25 79.945 57.313 ;
        RECT 72.606 47.636 72.652 64.606 ;
        RECT 55.638 64.604 72.606 64.652 ;
        RECT 63.038 57.204 79.991 57.267 ;
        RECT 72.56 47.682 72.606 64.652 ;
        RECT 55.592 64.65 72.56 64.698 ;
        RECT 63.084 57.158 80.037 57.221 ;
        RECT 72.514 47.728 72.56 64.698 ;
        RECT 55.546 64.696 72.514 64.744 ;
        RECT 63.13 57.112 80.083 57.175 ;
        RECT 72.468 47.774 72.514 64.744 ;
        RECT 55.5 64.742 72.468 64.79 ;
        RECT 63.176 57.066 80.129 57.129 ;
        RECT 72.422 47.82 72.468 64.79 ;
        RECT 55.454 64.788 72.422 64.836 ;
        RECT 63.222 57.02 80.175 57.083 ;
        RECT 72.376 47.866 72.422 64.836 ;
        RECT 55.408 64.834 72.376 64.882 ;
        RECT 63.268 56.974 80.221 57.037 ;
        RECT 72.33 47.912 72.376 64.882 ;
        RECT 55.362 64.88 72.33 64.928 ;
        RECT 63.314 56.928 80.267 56.991 ;
        RECT 72.284 47.958 72.33 64.928 ;
        RECT 55.316 64.926 72.284 64.974 ;
        RECT 63.36 56.882 80.313 56.945 ;
        RECT 72.238 48.004 72.284 64.974 ;
        RECT 55.27 64.972 72.238 65.02 ;
        RECT 63.406 56.836 80.359 56.899 ;
        RECT 72.192 48.05 72.238 65.02 ;
        RECT 55.224 65.018 72.192 65.066 ;
        RECT 63.452 56.79 80.405 56.853 ;
        RECT 72.146 48.096 72.192 65.066 ;
        RECT 55.178 65.064 72.146 65.112 ;
        RECT 63.498 56.744 80.451 56.807 ;
        RECT 72.1 48.142 72.146 65.112 ;
        RECT 55.132 65.11 72.1 65.158 ;
        RECT 63.544 56.698 80.497 56.761 ;
        RECT 72.054 48.188 72.1 65.158 ;
        RECT 55.086 65.156 72.054 65.204 ;
        RECT 63.59 56.652 80.543 56.715 ;
        RECT 72.008 48.234 72.054 65.204 ;
        RECT 55.04 65.202 72.008 65.25 ;
        RECT 63.636 56.606 80.589 56.669 ;
        RECT 71.962 48.28 72.008 65.25 ;
        RECT 54.994 65.248 71.962 65.296 ;
        RECT 63.682 56.56 80.635 56.623 ;
        RECT 71.916 48.326 71.962 65.296 ;
        RECT 54.948 65.294 71.916 65.342 ;
        RECT 63.728 56.514 80.681 56.577 ;
        RECT 71.87 48.372 71.916 65.342 ;
        RECT 54.902 65.34 71.87 65.388 ;
        RECT 63.774 56.468 80.727 56.531 ;
        RECT 71.824 48.418 71.87 65.388 ;
        RECT 54.856 65.386 71.824 65.434 ;
        RECT 63.82 56.422 80.773 56.485 ;
        RECT 71.778 48.464 71.824 65.434 ;
        RECT 54.81 65.432 71.778 65.48 ;
        RECT 63.866 56.376 80.819 56.439 ;
        RECT 71.732 48.51 71.778 65.48 ;
        RECT 54.764 65.478 71.732 65.526 ;
        RECT 63.912 56.33 80.865 56.393 ;
        RECT 71.686 48.556 71.732 65.526 ;
        RECT 54.718 65.524 71.686 65.572 ;
        RECT 63.958 56.284 80.911 56.347 ;
        RECT 71.64 48.602 71.686 65.572 ;
        RECT 54.672 65.57 71.64 65.618 ;
        RECT 64.004 56.238 80.957 56.301 ;
        RECT 71.594 48.648 71.64 65.618 ;
        RECT 54.626 65.616 71.594 65.664 ;
        RECT 64.05 56.192 81.003 56.255 ;
        RECT 71.548 48.694 71.594 65.664 ;
        RECT 54.58 65.662 71.548 65.71 ;
        RECT 64.096 56.146 81.049 56.209 ;
        RECT 71.502 48.74 71.548 65.71 ;
        RECT 54.534 65.708 71.502 65.756 ;
        RECT 64.142 56.1 81.095 56.163 ;
        RECT 71.456 48.786 71.502 65.756 ;
        RECT 54.488 65.754 71.456 65.802 ;
        RECT 64.188 56.054 81.141 56.117 ;
        RECT 71.41 48.832 71.456 65.802 ;
        RECT 54.442 65.8 71.41 65.848 ;
        RECT 64.234 56.008 81.187 56.071 ;
        RECT 71.364 48.878 71.41 65.848 ;
        RECT 54.396 65.846 71.364 65.894 ;
        RECT 64.28 55.962 81.233 56.024 ;
        RECT 71.318 48.924 71.364 65.894 ;
        RECT 54.35 65.892 71.318 65.94 ;
        RECT 64.326 55.916 110 56 ;
        RECT 71.272 48.97 71.318 65.94 ;
        RECT 54.304 65.938 71.272 65.986 ;
        RECT 64.372 55.87 110 56 ;
        RECT 71.226 49.016 71.272 65.986 ;
        RECT 54.258 65.984 71.226 66.032 ;
        RECT 64.418 55.824 110 56 ;
        RECT 71.18 49.062 71.226 66.032 ;
        RECT 54.212 66.03 71.18 66.078 ;
        RECT 64.464 55.778 110 56 ;
        RECT 71.134 49.108 71.18 66.078 ;
        RECT 54.166 66.076 71.134 66.124 ;
        RECT 64.51 55.732 110 56 ;
        RECT 71.088 49.154 71.134 66.124 ;
        RECT 54.12 66.122 71.088 66.17 ;
        RECT 64.556 55.686 110 56 ;
        RECT 71.042 49.2 71.088 66.17 ;
        RECT 54.074 66.168 71.042 66.216 ;
        RECT 64.602 55.64 110 56 ;
        RECT 70.996 49.246 71.042 66.216 ;
        RECT 54.028 66.214 70.996 66.262 ;
        RECT 64.648 55.594 110 56 ;
        RECT 70.95 49.292 70.996 66.262 ;
        RECT 53.982 66.26 70.95 66.308 ;
        RECT 64.694 55.548 110 56 ;
        RECT 70.904 49.338 70.95 66.308 ;
        RECT 53.936 66.306 70.904 66.354 ;
        RECT 64.74 55.502 110 56 ;
        RECT 70.858 49.384 70.904 66.354 ;
        RECT 53.89 66.352 70.858 66.4 ;
        RECT 64.786 55.456 110 56 ;
        RECT 70.812 49.43 70.858 66.4 ;
        RECT 53.844 66.398 70.812 66.446 ;
        RECT 64.832 55.41 110 56 ;
        RECT 70.766 49.476 70.812 66.446 ;
        RECT 53.798 66.444 70.766 66.492 ;
        RECT 64.878 55.364 110 56 ;
        RECT 70.72 49.522 70.766 66.492 ;
        RECT 53.752 66.49 70.72 66.538 ;
        RECT 64.924 55.318 110 56 ;
        RECT 70.674 49.568 70.72 66.538 ;
        RECT 53.706 66.536 70.674 66.584 ;
        RECT 64.97 55.272 110 56 ;
        RECT 70.628 49.614 70.674 66.584 ;
        RECT 53.66 66.582 70.628 66.63 ;
        RECT 65.016 55.226 110 56 ;
        RECT 70.582 49.66 70.628 66.63 ;
        RECT 53.614 66.628 70.582 66.676 ;
        RECT 65.062 55.18 110 56 ;
        RECT 70.536 49.706 70.582 66.676 ;
        RECT 53.568 66.674 70.536 66.722 ;
        RECT 65.108 55.134 110 56 ;
        RECT 70.49 49.752 70.536 66.722 ;
        RECT 53.522 66.72 70.49 66.768 ;
        RECT 65.154 55.088 110 56 ;
        RECT 70.444 49.798 70.49 66.768 ;
        RECT 53.476 66.766 70.444 66.814 ;
        RECT 65.2 55.042 110 56 ;
        RECT 70.398 49.844 70.444 66.814 ;
        RECT 53.43 66.812 70.398 66.86 ;
        RECT 65.246 54.996 110 56 ;
        RECT 70.352 49.89 70.398 66.86 ;
        RECT 53.384 66.858 70.352 66.906 ;
        RECT 65.292 54.95 110 56 ;
        RECT 70.306 49.936 70.352 66.906 ;
        RECT 53.338 66.904 70.306 66.952 ;
        RECT 65.338 54.904 110 56 ;
        RECT 70.26 49.982 70.306 66.952 ;
        RECT 53.292 66.95 70.26 66.998 ;
        RECT 65.384 54.858 110 56 ;
        RECT 70.214 50.028 70.26 66.998 ;
        RECT 53.246 66.996 70.214 67.044 ;
        RECT 65.43 54.812 110 56 ;
        RECT 70.168 50.074 70.214 67.044 ;
        RECT 53.2 67.042 70.168 67.09 ;
        RECT 65.476 54.766 110 56 ;
        RECT 70.122 50.12 70.168 67.09 ;
        RECT 53.154 67.088 70.122 67.136 ;
        RECT 65.522 54.72 110 56 ;
        RECT 70.076 50.166 70.122 67.136 ;
        RECT 53.108 67.134 70.076 67.182 ;
        RECT 65.568 54.674 110 56 ;
        RECT 70.03 50.212 70.076 67.182 ;
        RECT 53.062 67.18 70.03 67.228 ;
        RECT 65.614 54.628 110 56 ;
        RECT 69.984 50.258 70.03 67.228 ;
        RECT 53.016 67.226 69.984 67.274 ;
        RECT 65.66 54.582 110 56 ;
        RECT 69.938 50.304 69.984 67.274 ;
        RECT 52.97 67.272 69.938 67.32 ;
        RECT 65.706 54.536 110 56 ;
        RECT 69.892 50.35 69.938 67.32 ;
        RECT 52.924 67.318 69.892 67.366 ;
        RECT 65.752 54.49 110 56 ;
        RECT 69.846 50.396 69.892 67.366 ;
        RECT 52.878 67.364 69.846 67.412 ;
        RECT 65.798 54.444 110 56 ;
        RECT 69.8 50.442 69.846 67.412 ;
        RECT 52.832 67.41 69.8 67.458 ;
        RECT 65.844 54.398 110 56 ;
        RECT 69.754 50.488 69.8 67.458 ;
        RECT 52.786 67.456 69.754 67.504 ;
        RECT 65.89 54.352 110 56 ;
        RECT 69.708 50.534 69.754 67.504 ;
        RECT 52.74 67.502 69.708 67.55 ;
        RECT 65.936 54.306 110 56 ;
        RECT 69.662 50.58 69.708 67.55 ;
        RECT 52.694 67.548 69.662 67.596 ;
        RECT 65.982 54.26 110 56 ;
        RECT 69.616 50.626 69.662 67.596 ;
        RECT 52.648 67.594 69.616 67.642 ;
        RECT 66.028 54.214 110 56 ;
        RECT 69.57 50.672 69.616 67.642 ;
        RECT 52.602 67.64 69.57 67.688 ;
        RECT 66.074 54.168 110 56 ;
        RECT 69.524 50.718 69.57 67.688 ;
        RECT 52.556 67.686 69.524 67.734 ;
        RECT 66.12 54.122 110 56 ;
        RECT 69.478 50.764 69.524 67.734 ;
        RECT 52.51 67.732 69.478 67.78 ;
        RECT 66.166 54.076 110 56 ;
        RECT 69.432 50.81 69.478 67.78 ;
        RECT 52.464 67.778 69.432 67.826 ;
        RECT 66.212 54.03 110 56 ;
        RECT 69.386 50.856 69.432 67.826 ;
        RECT 52.418 67.824 69.386 67.872 ;
        RECT 66.258 53.984 110 56 ;
        RECT 69.34 50.902 69.386 67.872 ;
        RECT 52.372 67.87 69.34 67.918 ;
        RECT 66.304 53.938 110 56 ;
        RECT 69.294 50.948 69.34 67.918 ;
        RECT 52.326 67.916 69.294 67.964 ;
        RECT 66.35 53.892 110 56 ;
        RECT 69.248 50.994 69.294 67.964 ;
        RECT 52.28 67.962 69.248 68.01 ;
        RECT 66.396 53.846 110 56 ;
        RECT 69.202 51.04 69.248 68.01 ;
        RECT 52.234 68.008 69.202 68.056 ;
        RECT 66.442 53.8 110 56 ;
        RECT 69.156 51.086 69.202 68.056 ;
        RECT 52.188 68.054 69.156 68.102 ;
        RECT 66.488 53.754 110 56 ;
        RECT 69.11 51.132 69.156 68.102 ;
        RECT 52.142 68.1 69.11 68.148 ;
        RECT 66.534 53.708 110 56 ;
        RECT 69.064 51.178 69.11 68.148 ;
        RECT 52.096 68.146 69.064 68.194 ;
        RECT 66.58 53.662 110 56 ;
        RECT 69.018 51.224 69.064 68.194 ;
        RECT 52.05 68.192 69.018 68.24 ;
        RECT 66.626 53.616 110 56 ;
        RECT 68.972 51.27 69.018 68.24 ;
        RECT 52.004 68.238 68.972 68.286 ;
        RECT 66.672 53.57 110 56 ;
        RECT 68.926 51.316 68.972 68.286 ;
        RECT 51.958 68.284 68.926 68.332 ;
        RECT 66.718 53.524 110 56 ;
        RECT 68.88 51.362 68.926 68.332 ;
        RECT 51.912 68.33 68.88 68.378 ;
        RECT 66.764 53.478 110 56 ;
        RECT 68.834 51.408 68.88 68.378 ;
        RECT 51.866 68.376 68.834 68.424 ;
        RECT 66.81 53.432 110 56 ;
        RECT 68.788 51.454 68.834 68.424 ;
        RECT 51.82 68.422 68.788 68.47 ;
        RECT 66.856 53.386 110 56 ;
        RECT 68.742 51.5 68.788 68.47 ;
        RECT 51.774 68.468 68.742 68.516 ;
        RECT 66.902 53.34 110 56 ;
        RECT 68.696 51.546 68.742 68.516 ;
        RECT 51.728 68.514 68.696 68.562 ;
        RECT 66.948 53.294 110 56 ;
        RECT 68.65 51.592 68.696 68.562 ;
        RECT 51.682 68.56 68.65 68.608 ;
        RECT 66.994 53.248 110 56 ;
        RECT 68.604 51.638 68.65 68.608 ;
        RECT 51.636 68.606 68.604 68.654 ;
        RECT 67.04 53.202 110 56 ;
        RECT 68.558 51.684 68.604 68.654 ;
        RECT 51.59 68.652 68.558 68.7 ;
        RECT 67.086 53.156 110 56 ;
        RECT 68.512 51.73 68.558 68.7 ;
        RECT 51.544 68.698 68.512 68.746 ;
        RECT 67.132 53.11 110 56 ;
        RECT 68.466 51.776 68.512 68.746 ;
        RECT 51.498 68.744 68.466 68.792 ;
        RECT 67.178 53.064 110 56 ;
        RECT 68.42 51.822 68.466 68.792 ;
        RECT 51.452 68.79 68.42 68.838 ;
        RECT 67.224 53.018 110 56 ;
        RECT 68.374 51.868 68.42 68.838 ;
        RECT 51.406 68.836 68.374 68.884 ;
        RECT 67.27 52.972 110 56 ;
        RECT 68.328 51.914 68.374 68.884 ;
        RECT 51.36 68.882 68.328 68.93 ;
        RECT 67.316 52.926 110 56 ;
        RECT 68.282 51.96 68.328 68.93 ;
        RECT 51.314 68.928 68.282 68.976 ;
        RECT 67.362 52.88 110 56 ;
        RECT 68.236 52.006 68.282 68.976 ;
        RECT 51.268 68.974 68.236 69.022 ;
        RECT 67.408 52.834 110 56 ;
        RECT 68.19 52.052 68.236 69.022 ;
        RECT 51.222 69.02 68.19 69.068 ;
        RECT 67.454 52.788 110 56 ;
        RECT 68.144 52.098 68.19 69.068 ;
        RECT 51.176 69.066 68.144 69.114 ;
        RECT 67.5 52.742 110 56 ;
        RECT 68.098 52.144 68.144 69.114 ;
        RECT 51.13 69.112 68.098 69.16 ;
        RECT 67.546 52.696 110 56 ;
        RECT 68.052 52.19 68.098 69.16 ;
        RECT 51.084 69.158 68.052 69.206 ;
        RECT 67.592 52.65 110 56 ;
        RECT 68.006 52.236 68.052 69.206 ;
        RECT 51.038 69.204 68.006 69.252 ;
        RECT 67.638 52.604 110 56 ;
        RECT 67.96 52.282 68.006 69.252 ;
        RECT 50.992 69.25 67.96 69.298 ;
        RECT 67.684 52.558 110 56 ;
        RECT 67.914 52.328 67.96 69.298 ;
        RECT 50.946 69.296 67.914 69.344 ;
        RECT 67.73 52.512 110 56 ;
        RECT 67.868 52.374 67.914 69.344 ;
        RECT 50.9 69.342 67.868 69.39 ;
        RECT 67.776 52.466 110 56 ;
        RECT 67.822 52.42 67.868 69.39 ;
        RECT 50.854 69.388 67.822 69.436 ;
        RECT 50.808 69.434 67.776 69.482 ;
        RECT 50.762 69.48 67.73 69.528 ;
        RECT 50.716 69.526 67.684 69.574 ;
        RECT 50.67 69.572 67.638 69.62 ;
        RECT 50.624 69.618 67.592 69.666 ;
        RECT 50.578 69.664 67.546 69.712 ;
        RECT 50.532 69.71 67.5 69.758 ;
        RECT 50.486 69.756 67.454 69.804 ;
        RECT 50.44 69.802 67.408 69.85 ;
        RECT 50.394 69.848 67.362 69.896 ;
        RECT 50.348 69.894 67.316 69.942 ;
        RECT 50.302 69.94 67.27 69.988 ;
        RECT 50.256 69.986 67.224 70.034 ;
        RECT 50.21 70.032 67.178 70.08 ;
        RECT 50.164 70.078 67.132 70.126 ;
        RECT 50.118 70.124 67.086 70.172 ;
        RECT 50.072 70.17 67.04 70.218 ;
        RECT 50.026 70.216 66.994 70.264 ;
        RECT 49.98 70.262 66.948 70.31 ;
        RECT 49.934 70.308 66.902 70.356 ;
        RECT 49.888 70.354 66.856 70.402 ;
        RECT 49.842 70.4 66.81 70.448 ;
        RECT 49.796 70.446 66.764 70.494 ;
        RECT 49.75 70.492 66.718 70.54 ;
        RECT 49.704 70.538 66.672 70.586 ;
        RECT 49.658 70.584 66.626 70.632 ;
        RECT 49.612 70.63 66.58 70.678 ;
        RECT 49.566 70.676 66.534 70.724 ;
        RECT 49.52 70.722 66.488 70.77 ;
        RECT 49.474 70.768 66.442 70.816 ;
        RECT 49.428 70.814 66.396 70.862 ;
        RECT 49.382 70.86 66.35 70.908 ;
        RECT 49.336 70.906 66.304 70.954 ;
        RECT 49.29 70.952 66.258 71 ;
        RECT 49.244 70.998 66.212 71.046 ;
        RECT 49.198 71.044 66.166 71.092 ;
        RECT 49.152 71.09 66.12 71.138 ;
        RECT 49.106 71.136 66.074 71.184 ;
        RECT 49.06 71.182 66.028 71.23 ;
        RECT 49.014 71.228 65.982 71.276 ;
        RECT 48.968 71.274 65.936 71.322 ;
        RECT 48.922 71.32 65.89 71.368 ;
        RECT 48.876 71.366 65.844 71.414 ;
        RECT 48.83 71.412 65.798 71.46 ;
        RECT 48.784 71.458 65.752 71.506 ;
        RECT 48.738 71.504 65.706 71.552 ;
        RECT 48.692 71.55 65.66 71.598 ;
        RECT 48.646 71.596 65.614 71.644 ;
        RECT 48.6 71.642 65.568 71.69 ;
        RECT 48.554 71.688 65.522 71.736 ;
        RECT 48.508 71.734 65.476 71.782 ;
        RECT 48.462 71.78 65.43 71.828 ;
        RECT 48.416 71.826 65.384 71.874 ;
        RECT 48.37 71.872 65.338 71.92 ;
        RECT 48.324 71.918 65.292 71.966 ;
        RECT 48.278 71.964 65.246 72.012 ;
        RECT 48.232 72.01 65.2 72.058 ;
        RECT 48.186 72.056 65.154 72.104 ;
        RECT 48.14 72.102 65.108 72.15 ;
        RECT 48.094 72.148 65.062 72.196 ;
        RECT 48.048 72.194 65.016 72.242 ;
        RECT 48.002 72.24 64.97 72.288 ;
        RECT 47.956 72.286 64.924 72.334 ;
        RECT 47.91 72.332 64.878 72.38 ;
        RECT 47.864 72.378 64.832 72.426 ;
        RECT 47.818 72.424 64.786 72.472 ;
        RECT 47.772 72.47 64.74 72.518 ;
        RECT 47.726 72.516 64.694 72.564 ;
        RECT 47.68 72.562 64.648 72.61 ;
        RECT 47.634 72.608 64.602 72.656 ;
        RECT 47.588 72.654 64.556 72.702 ;
        RECT 47.542 72.7 64.51 72.748 ;
        RECT 47.496 72.746 64.464 72.794 ;
        RECT 47.45 72.792 64.418 72.84 ;
        RECT 47.404 72.838 64.372 72.886 ;
        RECT 47.358 72.884 64.326 72.932 ;
        RECT 47.312 72.93 64.28 72.978 ;
        RECT 47.266 72.976 64.234 73.024 ;
        RECT 47.22 73.022 64.188 73.07 ;
        RECT 47.174 73.068 64.142 73.116 ;
        RECT 47.128 73.114 64.096 73.162 ;
        RECT 47.082 73.16 64.05 73.208 ;
        RECT 47.036 73.206 64.004 73.254 ;
        RECT 46.99 73.252 63.958 73.3 ;
        RECT 46.944 73.298 63.912 73.346 ;
        RECT 46.898 73.344 63.866 73.392 ;
        RECT 46.852 73.39 63.82 73.438 ;
        RECT 46.806 73.436 63.774 73.484 ;
        RECT 46.76 73.482 63.728 73.53 ;
        RECT 46.714 73.528 63.682 73.576 ;
        RECT 46.668 73.574 63.636 73.622 ;
        RECT 46.622 73.62 63.59 73.668 ;
        RECT 46.576 73.666 63.544 73.714 ;
        RECT 46.53 73.712 63.498 73.76 ;
        RECT 46.484 73.758 63.452 73.806 ;
        RECT 46.438 73.804 63.406 73.852 ;
        RECT 46.392 73.85 63.36 73.898 ;
        RECT 46.346 73.896 63.314 73.944 ;
        RECT 46.3 73.942 63.268 73.99 ;
        RECT 46.254 73.988 63.222 74.036 ;
        RECT 46.208 74.034 63.176 74.082 ;
        RECT 46.162 74.08 63.13 74.128 ;
        RECT 46.116 74.126 63.084 74.174 ;
        RECT 46.07 74.172 63.038 74.22 ;
        RECT 46.024 74.218 62.992 74.266 ;
        RECT 45.978 74.264 62.946 74.312 ;
        RECT 45.932 74.31 62.9 74.358 ;
        RECT 45.886 74.356 62.854 74.404 ;
        RECT 45.84 74.402 62.808 74.45 ;
        RECT 45.794 74.448 62.762 74.496 ;
        RECT 45.748 74.494 62.716 74.542 ;
        RECT 45.702 74.54 62.67 74.588 ;
        RECT 45.656 74.586 62.624 74.634 ;
        RECT 45.61 74.632 62.578 74.68 ;
        RECT 45.564 74.678 62.532 74.726 ;
        RECT 45.518 74.724 62.486 74.772 ;
        RECT 45.472 74.77 62.44 74.818 ;
        RECT 45.426 74.816 62.394 74.864 ;
        RECT 45.38 74.862 62.348 74.91 ;
        RECT 45.334 74.908 62.302 74.956 ;
        RECT 45.288 74.954 62.256 75.002 ;
        RECT 45.242 75 62.21 75.048 ;
        RECT 45.196 75.046 62.164 75.094 ;
        RECT 45.15 75.092 62.118 75.14 ;
        RECT 45.104 75.138 62.072 75.186 ;
        RECT 45.058 75.184 62.026 75.232 ;
        RECT 45.012 75.23 61.98 75.278 ;
        RECT 44.966 75.276 61.934 75.324 ;
        RECT 44.92 75.322 61.888 75.37 ;
        RECT 44.874 75.368 61.842 75.416 ;
        RECT 44.828 75.414 61.796 75.462 ;
        RECT 44.782 75.46 61.75 75.508 ;
        RECT 44.736 75.506 61.704 75.554 ;
        RECT 44.69 75.552 61.658 75.6 ;
        RECT 44.644 75.598 61.612 75.646 ;
        RECT 44.598 75.644 61.566 75.692 ;
        RECT 44.552 75.69 61.52 75.738 ;
        RECT 44.506 75.736 61.474 75.784 ;
        RECT 44.46 75.782 61.428 75.83 ;
        RECT 44.414 75.828 61.382 75.876 ;
        RECT 44.368 75.874 61.336 75.922 ;
        RECT 44.322 75.92 61.29 75.968 ;
        RECT 44.276 75.966 61.244 76.014 ;
        RECT 44.23 76.012 61.198 76.06 ;
        RECT 44.184 76.058 61.152 76.106 ;
        RECT 44.138 76.104 61.106 76.152 ;
        RECT 44.092 76.15 61.06 76.198 ;
        RECT 44.046 76.196 61.014 76.244 ;
        RECT 44 76.242 60.968 76.29 ;
        RECT 44 76.242 60.922 76.336 ;
        RECT 44 76.242 60.876 76.382 ;
        RECT 44 76.242 60.83 76.428 ;
        RECT 44 76.242 60.784 76.474 ;
        RECT 44 76.242 60.738 76.52 ;
        RECT 44 76.242 60.692 76.566 ;
        RECT 44 76.242 60.646 76.612 ;
        RECT 44 76.242 60.6 76.658 ;
        RECT 44 76.242 60.554 76.704 ;
        RECT 44 76.242 60.508 76.75 ;
        RECT 44 76.242 60.462 76.796 ;
        RECT 44 76.242 60.416 76.842 ;
        RECT 44 76.242 60.37 76.888 ;
        RECT 44 76.242 60.324 76.934 ;
        RECT 44 76.242 60.278 76.98 ;
        RECT 44 76.242 60.232 77.026 ;
        RECT 44 76.242 60.186 77.072 ;
        RECT 44 76.242 60.14 77.118 ;
        RECT 44 76.242 60.094 77.164 ;
        RECT 44 76.242 60.048 77.21 ;
        RECT 44 76.242 60.002 77.256 ;
        RECT 44 76.242 59.956 77.302 ;
        RECT 44 76.242 59.91 77.348 ;
        RECT 44 76.242 59.864 77.394 ;
        RECT 44 76.242 59.818 77.44 ;
        RECT 44 76.242 59.772 77.486 ;
        RECT 44 76.242 59.726 77.532 ;
        RECT 44 76.242 59.68 77.578 ;
        RECT 44 76.242 59.634 77.624 ;
        RECT 44 76.242 59.588 77.67 ;
        RECT 44 76.242 59.542 77.716 ;
        RECT 44 76.242 59.496 77.762 ;
        RECT 44 76.242 59.45 77.808 ;
        RECT 44 76.242 59.404 77.854 ;
        RECT 44 76.242 59.358 77.9 ;
        RECT 44 76.242 59.312 77.946 ;
        RECT 44 76.242 59.266 77.992 ;
        RECT 44 76.242 59.22 78.038 ;
        RECT 44 76.242 59.174 78.084 ;
        RECT 44 76.242 59.128 78.13 ;
        RECT 44 76.242 59.082 78.176 ;
        RECT 44 76.242 59.036 78.222 ;
        RECT 44 76.242 58.99 78.268 ;
        RECT 44 76.242 58.944 78.314 ;
        RECT 44 76.242 58.898 78.36 ;
        RECT 44 76.242 58.852 78.406 ;
        RECT 44 76.242 58.806 78.452 ;
        RECT 44 76.242 58.76 78.498 ;
        RECT 44 76.242 58.714 78.544 ;
        RECT 44 76.242 58.668 78.59 ;
        RECT 44 76.242 58.622 78.636 ;
        RECT 44 76.242 58.576 78.682 ;
        RECT 44 76.242 58.53 78.728 ;
        RECT 44 76.242 58.484 78.774 ;
        RECT 44 76.242 58.438 78.82 ;
        RECT 44 76.242 58.392 78.866 ;
        RECT 44 76.242 58.346 78.912 ;
        RECT 44 76.242 58.3 78.958 ;
        RECT 44 76.242 58.254 79.004 ;
        RECT 44 76.242 58.208 79.05 ;
        RECT 44 76.242 58.162 79.096 ;
        RECT 44 76.242 58.116 79.142 ;
        RECT 44 76.242 58.07 79.188 ;
        RECT 44 76.242 58.024 79.234 ;
        RECT 44 76.242 57.978 79.28 ;
        RECT 44 76.242 57.932 79.326 ;
        RECT 44 76.242 57.886 79.372 ;
        RECT 44 76.242 57.84 79.418 ;
        RECT 44 76.242 57.794 79.464 ;
        RECT 44 76.242 57.748 79.51 ;
        RECT 44 76.242 57.702 79.556 ;
        RECT 44 76.242 57.656 79.602 ;
        RECT 44 76.242 57.61 79.648 ;
        RECT 44 76.242 57.564 79.694 ;
        RECT 44 76.242 57.518 79.74 ;
        RECT 44 76.242 57.472 79.786 ;
        RECT 44 76.242 57.426 79.832 ;
        RECT 44 76.242 57.38 79.878 ;
        RECT 44 76.242 57.334 79.924 ;
        RECT 44 76.242 57.288 79.97 ;
        RECT 44 76.242 57.242 80.016 ;
        RECT 44 76.242 57.196 80.062 ;
        RECT 44 76.242 57.15 80.108 ;
        RECT 44 76.242 57.104 80.154 ;
        RECT 44 76.242 57.058 80.2 ;
        RECT 44 76.242 57.012 80.246 ;
        RECT 44 76.242 56.966 80.292 ;
        RECT 44 76.242 56.92 80.338 ;
        RECT 44 76.242 56.874 80.384 ;
        RECT 44 76.242 56.828 80.43 ;
        RECT 44 76.242 56.782 80.476 ;
        RECT 44 76.242 56.736 80.522 ;
        RECT 44 76.242 56.69 80.568 ;
        RECT 44 76.242 56.644 80.614 ;
        RECT 44 76.242 56.598 80.66 ;
        RECT 44 76.242 56.552 80.706 ;
        RECT 44 76.242 56.506 80.752 ;
        RECT 44 76.242 56.46 80.798 ;
        RECT 44 76.242 56.414 80.844 ;
        RECT 44 76.242 56.368 80.89 ;
        RECT 44 76.242 56.322 80.936 ;
        RECT 44 76.242 56.276 80.982 ;
        RECT 44 76.242 56.23 81.028 ;
        RECT 44 76.242 56.184 81.074 ;
        RECT 44 76.242 56.138 81.12 ;
        RECT 44 76.242 56.092 81.166 ;
        RECT 44 76.242 56.046 81.212 ;
        RECT 44 76.242 56 110 ;
        RECT 82.76 57.5 110 63.5 ;
        RECT 76.748 63.489 85.24 63.521 ;
        RECT 74.31 65.927 82.76 65.996 ;
        RECT 74.356 65.881 82.806 65.957 ;
        RECT 82.728 57.516 82.76 65.996 ;
        RECT 74.264 65.973 82.728 66.035 ;
        RECT 74.402 65.835 82.852 65.911 ;
        RECT 82.682 57.555 82.728 66.035 ;
        RECT 74.218 66.019 82.682 66.081 ;
        RECT 74.448 65.789 82.898 65.865 ;
        RECT 82.636 57.601 82.682 66.081 ;
        RECT 74.172 66.065 82.636 66.127 ;
        RECT 74.494 65.743 82.944 65.819 ;
        RECT 82.59 57.647 82.636 66.127 ;
        RECT 74.126 66.111 82.59 66.173 ;
        RECT 74.54 65.697 82.99 65.773 ;
        RECT 82.544 57.693 82.59 66.173 ;
        RECT 74.08 66.157 82.544 66.219 ;
        RECT 74.586 65.651 83.036 65.727 ;
        RECT 82.498 57.739 82.544 66.219 ;
        RECT 74.034 66.203 82.498 66.265 ;
        RECT 74.632 65.605 83.082 65.681 ;
        RECT 82.452 57.785 82.498 66.265 ;
        RECT 73.988 66.249 82.452 66.311 ;
        RECT 74.678 65.559 83.128 65.635 ;
        RECT 82.406 57.831 82.452 66.311 ;
        RECT 73.942 66.295 82.406 66.357 ;
        RECT 74.724 65.513 83.174 65.589 ;
        RECT 82.36 57.877 82.406 66.357 ;
        RECT 73.896 66.341 82.36 66.403 ;
        RECT 74.77 65.467 83.22 65.543 ;
        RECT 82.314 57.923 82.36 66.403 ;
        RECT 73.85 66.387 82.314 66.449 ;
        RECT 74.816 65.421 83.266 65.497 ;
        RECT 82.268 57.969 82.314 66.449 ;
        RECT 73.804 66.433 82.268 66.495 ;
        RECT 74.862 65.375 83.312 65.451 ;
        RECT 82.222 58.015 82.268 66.495 ;
        RECT 73.758 66.479 82.222 66.541 ;
        RECT 74.908 65.329 83.358 65.405 ;
        RECT 82.176 58.061 82.222 66.541 ;
        RECT 73.712 66.525 82.176 66.587 ;
        RECT 74.954 65.283 83.404 65.359 ;
        RECT 82.13 58.107 82.176 66.587 ;
        RECT 73.666 66.571 82.13 66.633 ;
        RECT 75 65.237 83.45 65.313 ;
        RECT 82.084 58.153 82.13 66.633 ;
        RECT 73.62 66.617 82.084 66.679 ;
        RECT 75.046 65.191 83.496 65.267 ;
        RECT 82.038 58.199 82.084 66.679 ;
        RECT 73.574 66.663 82.038 66.725 ;
        RECT 75.092 65.145 83.542 65.221 ;
        RECT 81.992 58.245 82.038 66.725 ;
        RECT 73.528 66.709 81.992 66.771 ;
        RECT 75.138 65.099 83.588 65.175 ;
        RECT 81.946 58.291 81.992 66.771 ;
        RECT 73.482 66.755 81.946 66.817 ;
        RECT 75.184 65.053 83.634 65.129 ;
        RECT 81.9 58.337 81.946 66.817 ;
        RECT 73.436 66.801 81.9 66.863 ;
        RECT 75.23 65.007 83.68 65.083 ;
        RECT 81.854 58.383 81.9 66.863 ;
        RECT 73.39 66.847 81.854 66.909 ;
        RECT 75.276 64.961 83.726 65.037 ;
        RECT 81.808 58.429 81.854 66.909 ;
        RECT 73.344 66.893 81.808 66.955 ;
        RECT 75.322 64.915 83.772 64.991 ;
        RECT 81.762 58.475 81.808 66.955 ;
        RECT 73.298 66.939 81.762 67.001 ;
        RECT 75.368 64.869 83.818 64.945 ;
        RECT 81.716 58.521 81.762 67.001 ;
        RECT 73.252 66.985 81.716 67.047 ;
        RECT 75.414 64.823 83.864 64.899 ;
        RECT 81.67 58.567 81.716 67.047 ;
        RECT 73.206 67.031 81.67 67.093 ;
        RECT 75.46 64.777 83.91 64.853 ;
        RECT 81.624 58.613 81.67 67.093 ;
        RECT 73.16 67.077 81.624 67.139 ;
        RECT 75.506 64.731 83.956 64.807 ;
        RECT 81.578 58.659 81.624 67.139 ;
        RECT 73.114 67.123 81.578 67.185 ;
        RECT 75.552 64.685 84.002 64.761 ;
        RECT 81.532 58.705 81.578 67.185 ;
        RECT 73.068 67.169 81.532 67.231 ;
        RECT 75.598 64.639 84.048 64.715 ;
        RECT 81.486 58.751 81.532 67.231 ;
        RECT 73.022 67.215 81.486 67.277 ;
        RECT 75.644 64.593 84.094 64.669 ;
        RECT 81.44 58.797 81.486 67.277 ;
        RECT 72.976 67.261 81.44 67.323 ;
        RECT 75.69 64.547 84.14 64.623 ;
        RECT 81.394 58.843 81.44 67.323 ;
        RECT 72.93 67.307 81.394 67.369 ;
        RECT 75.736 64.501 84.186 64.577 ;
        RECT 81.348 58.889 81.394 67.369 ;
        RECT 72.884 67.353 81.348 67.415 ;
        RECT 75.782 64.455 84.232 64.531 ;
        RECT 81.302 58.935 81.348 67.415 ;
        RECT 72.838 67.399 81.302 67.461 ;
        RECT 75.828 64.409 84.278 64.485 ;
        RECT 81.256 58.981 81.302 67.461 ;
        RECT 72.792 67.445 81.256 67.507 ;
        RECT 75.874 64.363 84.324 64.439 ;
        RECT 81.21 59.027 81.256 67.507 ;
        RECT 72.746 67.491 81.21 67.553 ;
        RECT 75.92 64.317 84.37 64.393 ;
        RECT 81.164 59.073 81.21 67.553 ;
        RECT 72.7 67.537 81.164 67.599 ;
        RECT 75.966 64.271 84.416 64.347 ;
        RECT 81.118 59.119 81.164 67.599 ;
        RECT 72.654 67.583 81.118 67.645 ;
        RECT 76.012 64.225 84.462 64.301 ;
        RECT 81.072 59.165 81.118 67.645 ;
        RECT 72.608 67.629 81.072 67.691 ;
        RECT 76.058 64.179 84.508 64.255 ;
        RECT 81.026 59.211 81.072 67.691 ;
        RECT 72.562 67.675 81.026 67.737 ;
        RECT 76.104 64.133 84.554 64.209 ;
        RECT 80.98 59.257 81.026 67.737 ;
        RECT 72.516 67.721 80.98 67.783 ;
        RECT 76.15 64.087 84.6 64.163 ;
        RECT 80.934 59.303 80.98 67.783 ;
        RECT 72.47 67.767 80.934 67.829 ;
        RECT 76.196 64.041 84.646 64.117 ;
        RECT 80.888 59.349 80.934 67.829 ;
        RECT 72.424 67.813 80.888 67.875 ;
        RECT 76.242 63.995 84.692 64.071 ;
        RECT 80.842 59.395 80.888 67.875 ;
        RECT 72.378 67.859 80.842 67.921 ;
        RECT 76.288 63.949 84.738 64.025 ;
        RECT 80.796 59.441 80.842 67.921 ;
        RECT 72.332 67.905 80.796 67.967 ;
        RECT 76.334 63.903 84.784 63.979 ;
        RECT 80.75 59.487 80.796 67.967 ;
        RECT 72.286 67.951 80.75 68.013 ;
        RECT 76.38 63.857 84.83 63.933 ;
        RECT 80.704 59.533 80.75 68.013 ;
        RECT 72.24 67.997 80.704 68.059 ;
        RECT 76.426 63.811 84.876 63.887 ;
        RECT 80.658 59.579 80.704 68.059 ;
        RECT 72.194 68.043 80.658 68.105 ;
        RECT 76.472 63.765 84.922 63.841 ;
        RECT 80.612 59.625 80.658 68.105 ;
        RECT 72.148 68.089 80.612 68.151 ;
        RECT 76.518 63.719 84.968 63.795 ;
        RECT 80.566 59.671 80.612 68.151 ;
        RECT 72.102 68.135 80.566 68.197 ;
        RECT 76.564 63.673 85.014 63.749 ;
        RECT 80.52 59.717 80.566 68.197 ;
        RECT 72.056 68.181 80.52 68.243 ;
        RECT 76.61 63.627 85.06 63.703 ;
        RECT 80.474 59.763 80.52 68.243 ;
        RECT 72.01 68.227 80.474 68.289 ;
        RECT 76.656 63.581 85.106 63.657 ;
        RECT 80.428 59.809 80.474 68.289 ;
        RECT 71.964 68.273 80.428 68.335 ;
        RECT 76.702 63.535 85.152 63.611 ;
        RECT 80.382 59.855 80.428 68.335 ;
        RECT 71.918 68.319 80.382 68.381 ;
        RECT 76.748 63.489 85.198 63.565 ;
        RECT 80.336 59.901 80.382 68.381 ;
        RECT 71.872 68.365 80.336 68.427 ;
        RECT 76.794 63.443 110 63.5 ;
        RECT 80.29 59.947 80.336 68.427 ;
        RECT 71.826 68.411 80.29 68.473 ;
        RECT 76.84 63.397 110 63.5 ;
        RECT 80.244 59.993 80.29 68.473 ;
        RECT 71.78 68.457 80.244 68.519 ;
        RECT 76.886 63.351 110 63.5 ;
        RECT 80.198 60.039 80.244 68.519 ;
        RECT 71.734 68.503 80.198 68.565 ;
        RECT 76.932 63.305 110 63.5 ;
        RECT 80.152 60.085 80.198 68.565 ;
        RECT 71.688 68.549 80.152 68.611 ;
        RECT 76.978 63.259 110 63.5 ;
        RECT 80.106 60.131 80.152 68.611 ;
        RECT 71.642 68.595 80.106 68.657 ;
        RECT 77.024 63.213 110 63.5 ;
        RECT 80.06 60.177 80.106 68.657 ;
        RECT 71.596 68.641 80.06 68.703 ;
        RECT 77.07 63.167 110 63.5 ;
        RECT 80.014 60.223 80.06 68.703 ;
        RECT 71.55 68.687 80.014 68.749 ;
        RECT 77.116 63.121 110 63.5 ;
        RECT 79.968 60.269 80.014 68.749 ;
        RECT 71.504 68.733 79.968 68.795 ;
        RECT 77.162 63.075 110 63.5 ;
        RECT 79.922 60.315 79.968 68.795 ;
        RECT 71.458 68.779 79.922 68.841 ;
        RECT 77.208 63.029 110 63.5 ;
        RECT 79.876 60.361 79.922 68.841 ;
        RECT 71.412 68.825 79.876 68.887 ;
        RECT 77.254 62.983 110 63.5 ;
        RECT 79.83 60.407 79.876 68.887 ;
        RECT 71.366 68.871 79.83 68.933 ;
        RECT 77.3 62.937 110 63.5 ;
        RECT 79.784 60.453 79.83 68.933 ;
        RECT 71.32 68.917 79.784 68.979 ;
        RECT 77.346 62.891 110 63.5 ;
        RECT 79.738 60.499 79.784 68.979 ;
        RECT 71.274 68.963 79.738 69.025 ;
        RECT 77.392 62.845 110 63.5 ;
        RECT 79.692 60.545 79.738 69.025 ;
        RECT 71.228 69.009 79.692 69.071 ;
        RECT 77.438 62.799 110 63.5 ;
        RECT 79.646 60.591 79.692 69.071 ;
        RECT 71.182 69.055 79.646 69.117 ;
        RECT 77.484 62.753 110 63.5 ;
        RECT 79.6 60.637 79.646 69.117 ;
        RECT 71.136 69.101 79.6 69.163 ;
        RECT 77.53 62.707 110 63.5 ;
        RECT 79.554 60.683 79.6 69.163 ;
        RECT 71.09 69.147 79.554 69.209 ;
        RECT 77.576 62.661 110 63.5 ;
        RECT 79.508 60.729 79.554 69.209 ;
        RECT 71.044 69.193 79.508 69.255 ;
        RECT 77.622 62.615 110 63.5 ;
        RECT 79.462 60.775 79.508 69.255 ;
        RECT 70.998 69.239 79.462 69.301 ;
        RECT 77.668 62.569 110 63.5 ;
        RECT 79.416 60.821 79.462 69.301 ;
        RECT 70.952 69.285 79.416 69.347 ;
        RECT 77.714 62.523 110 63.5 ;
        RECT 79.37 60.867 79.416 69.347 ;
        RECT 70.906 69.331 79.37 69.393 ;
        RECT 77.76 62.477 110 63.5 ;
        RECT 79.324 60.913 79.37 69.393 ;
        RECT 70.86 69.377 79.324 69.439 ;
        RECT 77.806 62.431 110 63.5 ;
        RECT 79.278 60.959 79.324 69.439 ;
        RECT 69.515 30.5 110 42.5 ;
        RECT 57.496 42.496 74.483 42.524 ;
        RECT 52.574 47.418 69.515 47.477 ;
        RECT 52.62 47.372 69.561 47.447 ;
        RECT 69.502 30.506 69.515 47.477 ;
        RECT 52.666 47.326 69.607 47.401 ;
        RECT 69.456 30.536 69.502 47.506 ;
        RECT 52.528 47.464 69.456 47.552 ;
        RECT 52.712 47.28 69.653 47.355 ;
        RECT 69.41 30.582 69.456 47.552 ;
        RECT 52.482 47.51 69.41 47.598 ;
        RECT 52.758 47.234 69.699 47.309 ;
        RECT 69.364 30.628 69.41 47.598 ;
        RECT 52.436 47.556 69.364 47.644 ;
        RECT 52.804 47.188 69.745 47.263 ;
        RECT 69.318 30.674 69.364 47.644 ;
        RECT 52.39 47.602 69.318 47.69 ;
        RECT 52.85 47.142 69.791 47.217 ;
        RECT 69.272 30.72 69.318 47.69 ;
        RECT 52.344 47.648 69.272 47.736 ;
        RECT 52.896 47.096 69.837 47.171 ;
        RECT 69.226 30.766 69.272 47.736 ;
        RECT 52.298 47.694 69.226 47.782 ;
        RECT 52.942 47.05 69.883 47.125 ;
        RECT 69.18 30.812 69.226 47.782 ;
        RECT 52.252 47.74 69.18 47.828 ;
        RECT 52.988 47.004 69.929 47.079 ;
        RECT 69.134 30.858 69.18 47.828 ;
        RECT 52.206 47.786 69.134 47.874 ;
        RECT 53.034 46.958 69.975 47.033 ;
        RECT 69.088 30.904 69.134 47.874 ;
        RECT 52.16 47.832 69.088 47.92 ;
        RECT 53.08 46.912 70.021 46.987 ;
        RECT 69.042 30.95 69.088 47.92 ;
        RECT 52.114 47.878 69.042 47.966 ;
        RECT 53.126 46.866 70.067 46.941 ;
        RECT 68.996 30.996 69.042 47.966 ;
        RECT 52.068 47.924 68.996 48.012 ;
        RECT 53.172 46.82 70.113 46.895 ;
        RECT 68.95 31.042 68.996 48.012 ;
        RECT 52.022 47.97 68.95 48.058 ;
        RECT 53.218 46.774 70.159 46.849 ;
        RECT 68.904 31.088 68.95 48.058 ;
        RECT 51.976 48.016 68.904 48.104 ;
        RECT 53.264 46.728 70.205 46.803 ;
        RECT 68.858 31.134 68.904 48.104 ;
        RECT 51.93 48.062 68.858 48.15 ;
        RECT 53.31 46.682 70.251 46.757 ;
        RECT 68.812 31.18 68.858 48.15 ;
        RECT 51.884 48.108 68.812 48.196 ;
        RECT 53.356 46.636 70.297 46.711 ;
        RECT 68.766 31.226 68.812 48.196 ;
        RECT 51.838 48.154 68.766 48.242 ;
        RECT 53.402 46.59 70.343 46.665 ;
        RECT 68.72 31.272 68.766 48.242 ;
        RECT 51.792 48.2 68.72 48.288 ;
        RECT 53.448 46.544 70.389 46.619 ;
        RECT 68.674 31.318 68.72 48.288 ;
        RECT 51.746 48.246 68.674 48.334 ;
        RECT 53.494 46.498 70.435 46.573 ;
        RECT 68.628 31.364 68.674 48.334 ;
        RECT 51.7 48.292 68.628 48.38 ;
        RECT 53.54 46.452 70.481 46.527 ;
        RECT 68.582 31.41 68.628 48.38 ;
        RECT 51.654 48.338 68.582 48.426 ;
        RECT 53.586 46.406 70.527 46.481 ;
        RECT 68.536 31.456 68.582 48.426 ;
        RECT 51.608 48.384 68.536 48.472 ;
        RECT 53.632 46.36 70.573 46.435 ;
        RECT 68.49 31.502 68.536 48.472 ;
        RECT 51.562 48.43 68.49 48.518 ;
        RECT 53.678 46.314 70.619 46.389 ;
        RECT 68.444 31.548 68.49 48.518 ;
        RECT 51.516 48.476 68.444 48.564 ;
        RECT 53.724 46.268 70.665 46.343 ;
        RECT 68.398 31.594 68.444 48.564 ;
        RECT 51.47 48.522 68.398 48.61 ;
        RECT 53.77 46.222 70.711 46.297 ;
        RECT 68.352 31.64 68.398 48.61 ;
        RECT 51.424 48.568 68.352 48.656 ;
        RECT 53.816 46.176 70.757 46.251 ;
        RECT 68.306 31.686 68.352 48.656 ;
        RECT 51.378 48.614 68.306 48.702 ;
        RECT 53.862 46.13 70.803 46.205 ;
        RECT 68.26 31.732 68.306 48.702 ;
        RECT 51.332 48.66 68.26 48.748 ;
        RECT 53.908 46.084 70.849 46.159 ;
        RECT 68.214 31.778 68.26 48.748 ;
        RECT 51.286 48.706 68.214 48.794 ;
        RECT 53.954 46.038 70.895 46.113 ;
        RECT 68.168 31.824 68.214 48.794 ;
        RECT 51.24 48.752 68.168 48.84 ;
        RECT 54 45.992 70.941 46.067 ;
        RECT 68.122 31.87 68.168 48.84 ;
        RECT 51.194 48.798 68.122 48.886 ;
        RECT 54.046 45.946 70.987 46.021 ;
        RECT 68.076 31.916 68.122 48.886 ;
        RECT 51.148 48.844 68.076 48.932 ;
        RECT 54.092 45.9 71.033 45.975 ;
        RECT 68.03 31.962 68.076 48.932 ;
        RECT 51.102 48.89 68.03 48.978 ;
        RECT 54.138 45.854 71.079 45.929 ;
        RECT 67.984 32.008 68.03 48.978 ;
        RECT 51.056 48.936 67.984 49.024 ;
        RECT 54.184 45.808 71.125 45.883 ;
        RECT 67.938 32.054 67.984 49.024 ;
        RECT 51.01 48.982 67.938 49.07 ;
        RECT 54.23 45.762 71.171 45.837 ;
        RECT 67.892 32.1 67.938 49.07 ;
        RECT 50.964 49.028 67.892 49.116 ;
        RECT 54.276 45.716 71.217 45.791 ;
        RECT 67.846 32.146 67.892 49.116 ;
        RECT 50.918 49.074 67.846 49.162 ;
        RECT 54.322 45.67 71.263 45.745 ;
        RECT 67.8 32.192 67.846 49.162 ;
        RECT 50.872 49.12 67.8 49.208 ;
        RECT 54.368 45.624 71.309 45.699 ;
        RECT 67.754 32.238 67.8 49.208 ;
        RECT 50.826 49.166 67.754 49.254 ;
        RECT 54.414 45.578 71.355 45.653 ;
        RECT 67.708 32.284 67.754 49.254 ;
        RECT 50.78 49.212 67.708 49.3 ;
        RECT 54.46 45.532 71.401 45.607 ;
        RECT 67.662 32.33 67.708 49.3 ;
        RECT 50.734 49.258 67.662 49.346 ;
        RECT 54.506 45.486 71.447 45.561 ;
        RECT 67.616 32.376 67.662 49.346 ;
        RECT 50.688 49.304 67.616 49.392 ;
        RECT 54.552 45.44 71.493 45.515 ;
        RECT 67.57 32.422 67.616 49.392 ;
        RECT 50.642 49.35 67.57 49.438 ;
        RECT 54.598 45.394 71.539 45.469 ;
        RECT 67.524 32.468 67.57 49.438 ;
        RECT 50.596 49.396 67.524 49.484 ;
        RECT 54.644 45.348 71.585 45.423 ;
        RECT 67.478 32.514 67.524 49.484 ;
        RECT 50.55 49.442 67.478 49.53 ;
        RECT 54.69 45.302 71.631 45.377 ;
        RECT 67.432 32.56 67.478 49.53 ;
        RECT 50.504 49.488 67.432 49.576 ;
        RECT 54.736 45.256 71.677 45.331 ;
        RECT 67.386 32.606 67.432 49.576 ;
        RECT 50.458 49.534 67.386 49.622 ;
        RECT 54.782 45.21 71.723 45.285 ;
        RECT 67.34 32.652 67.386 49.622 ;
        RECT 50.412 49.58 67.34 49.668 ;
        RECT 54.828 45.164 71.769 45.239 ;
        RECT 67.294 32.698 67.34 49.668 ;
        RECT 50.366 49.626 67.294 49.714 ;
        RECT 54.874 45.118 71.815 45.193 ;
        RECT 67.248 32.744 67.294 49.714 ;
        RECT 50.32 49.672 67.248 49.76 ;
        RECT 54.92 45.072 71.861 45.147 ;
        RECT 67.202 32.79 67.248 49.76 ;
        RECT 50.274 49.718 67.202 49.806 ;
        RECT 54.966 45.026 71.907 45.101 ;
        RECT 67.156 32.836 67.202 49.806 ;
        RECT 50.228 49.764 67.156 49.852 ;
        RECT 55.012 44.98 71.953 45.055 ;
        RECT 67.11 32.882 67.156 49.852 ;
        RECT 50.182 49.81 67.11 49.898 ;
        RECT 55.058 44.934 71.999 45.009 ;
        RECT 67.064 32.928 67.11 49.898 ;
        RECT 50.136 49.856 67.064 49.944 ;
        RECT 55.104 44.888 72.045 44.963 ;
        RECT 67.018 32.974 67.064 49.944 ;
        RECT 50.09 49.902 67.018 49.99 ;
        RECT 55.15 44.842 72.091 44.917 ;
        RECT 66.972 33.02 67.018 49.99 ;
        RECT 50.044 49.948 66.972 50.036 ;
        RECT 55.196 44.796 72.137 44.871 ;
        RECT 66.926 33.066 66.972 50.036 ;
        RECT 49.998 49.994 66.926 50.082 ;
        RECT 55.242 44.75 72.183 44.825 ;
        RECT 66.88 33.112 66.926 50.082 ;
        RECT 49.952 50.04 66.88 50.128 ;
        RECT 55.288 44.704 72.229 44.779 ;
        RECT 66.834 33.158 66.88 50.128 ;
        RECT 49.906 50.086 66.834 50.174 ;
        RECT 55.334 44.658 72.275 44.733 ;
        RECT 66.788 33.204 66.834 50.174 ;
        RECT 49.86 50.132 66.788 50.22 ;
        RECT 55.38 44.612 72.321 44.687 ;
        RECT 66.742 33.25 66.788 50.22 ;
        RECT 49.814 50.178 66.742 50.266 ;
        RECT 55.426 44.566 72.367 44.641 ;
        RECT 66.696 33.296 66.742 50.266 ;
        RECT 49.768 50.224 66.696 50.312 ;
        RECT 55.472 44.52 72.413 44.595 ;
        RECT 66.65 33.342 66.696 50.312 ;
        RECT 49.722 50.27 66.65 50.358 ;
        RECT 55.518 44.474 72.459 44.549 ;
        RECT 66.604 33.388 66.65 50.358 ;
        RECT 49.676 50.316 66.604 50.404 ;
        RECT 55.564 44.428 72.505 44.503 ;
        RECT 66.558 33.434 66.604 50.404 ;
        RECT 49.63 50.362 66.558 50.45 ;
        RECT 55.61 44.382 72.551 44.457 ;
        RECT 66.512 33.48 66.558 50.45 ;
        RECT 49.584 50.408 66.512 50.496 ;
        RECT 55.656 44.336 72.597 44.411 ;
        RECT 66.466 33.526 66.512 50.496 ;
        RECT 49.538 50.454 66.466 50.542 ;
        RECT 55.702 44.29 72.643 44.365 ;
        RECT 66.42 33.572 66.466 50.542 ;
        RECT 49.492 50.5 66.42 50.588 ;
        RECT 55.748 44.244 72.689 44.319 ;
        RECT 66.374 33.618 66.42 50.588 ;
        RECT 49.446 50.546 66.374 50.634 ;
        RECT 55.794 44.198 72.735 44.273 ;
        RECT 66.328 33.664 66.374 50.634 ;
        RECT 49.4 50.592 66.328 50.68 ;
        RECT 55.84 44.152 72.781 44.227 ;
        RECT 66.282 33.71 66.328 50.68 ;
        RECT 49.354 50.638 66.282 50.726 ;
        RECT 55.886 44.106 72.827 44.181 ;
        RECT 66.236 33.756 66.282 50.726 ;
        RECT 49.308 50.684 66.236 50.772 ;
        RECT 55.932 44.06 72.873 44.135 ;
        RECT 66.19 33.802 66.236 50.772 ;
        RECT 49.262 50.73 66.19 50.818 ;
        RECT 55.978 44.014 72.919 44.089 ;
        RECT 66.144 33.848 66.19 50.818 ;
        RECT 49.216 50.776 66.144 50.864 ;
        RECT 56.024 43.968 72.965 44.043 ;
        RECT 66.098 33.894 66.144 50.864 ;
        RECT 49.17 50.822 66.098 50.91 ;
        RECT 56.07 43.922 73.011 43.997 ;
        RECT 66.052 33.94 66.098 50.91 ;
        RECT 49.124 50.868 66.052 50.956 ;
        RECT 56.116 43.876 73.057 43.951 ;
        RECT 66.006 33.986 66.052 50.956 ;
        RECT 49.078 50.914 66.006 51.002 ;
        RECT 56.162 43.83 73.103 43.905 ;
        RECT 65.96 34.032 66.006 51.002 ;
        RECT 49.032 50.96 65.96 51.048 ;
        RECT 56.208 43.784 73.149 43.859 ;
        RECT 65.914 34.078 65.96 51.048 ;
        RECT 48.986 51.006 65.914 51.094 ;
        RECT 56.254 43.738 73.195 43.813 ;
        RECT 65.868 34.124 65.914 51.094 ;
        RECT 48.94 51.052 65.868 51.14 ;
        RECT 56.3 43.692 73.241 43.767 ;
        RECT 65.822 34.17 65.868 51.14 ;
        RECT 48.894 51.098 65.822 51.186 ;
        RECT 56.346 43.646 73.287 43.721 ;
        RECT 65.776 34.216 65.822 51.186 ;
        RECT 48.848 51.144 65.776 51.232 ;
        RECT 56.392 43.6 73.333 43.675 ;
        RECT 65.73 34.262 65.776 51.232 ;
        RECT 48.802 51.19 65.73 51.278 ;
        RECT 56.438 43.554 73.379 43.629 ;
        RECT 65.684 34.308 65.73 51.278 ;
        RECT 48.756 51.236 65.684 51.324 ;
        RECT 56.484 43.508 73.425 43.583 ;
        RECT 65.638 34.354 65.684 51.324 ;
        RECT 48.71 51.282 65.638 51.37 ;
        RECT 56.53 43.462 73.471 43.537 ;
        RECT 65.592 34.4 65.638 51.37 ;
        RECT 48.664 51.328 65.592 51.416 ;
        RECT 56.576 43.416 73.517 43.491 ;
        RECT 65.546 34.446 65.592 51.416 ;
        RECT 48.618 51.374 65.546 51.462 ;
        RECT 56.622 43.37 73.563 43.445 ;
        RECT 65.5 34.492 65.546 51.462 ;
        RECT 48.572 51.42 65.5 51.508 ;
        RECT 56.668 43.324 73.609 43.399 ;
        RECT 65.454 34.538 65.5 51.508 ;
        RECT 48.526 51.466 65.454 51.554 ;
        RECT 56.714 43.278 73.655 43.353 ;
        RECT 65.408 34.584 65.454 51.554 ;
        RECT 48.48 51.512 65.408 51.6 ;
        RECT 56.76 43.232 73.701 43.307 ;
        RECT 65.362 34.63 65.408 51.6 ;
        RECT 48.434 51.558 65.362 51.646 ;
        RECT 56.806 43.186 73.747 43.261 ;
        RECT 65.316 34.676 65.362 51.646 ;
        RECT 48.388 51.604 65.316 51.692 ;
        RECT 56.852 43.14 73.793 43.215 ;
        RECT 65.27 34.722 65.316 51.692 ;
        RECT 48.342 51.65 65.27 51.738 ;
        RECT 56.898 43.094 73.839 43.169 ;
        RECT 65.224 34.768 65.27 51.738 ;
        RECT 48.296 51.696 65.224 51.784 ;
        RECT 56.944 43.048 73.885 43.123 ;
        RECT 65.178 34.814 65.224 51.784 ;
        RECT 48.25 51.742 65.178 51.83 ;
        RECT 56.99 43.002 73.931 43.077 ;
        RECT 65.132 34.86 65.178 51.83 ;
        RECT 48.204 51.788 65.132 51.876 ;
        RECT 57.036 42.956 73.977 43.031 ;
        RECT 65.086 34.906 65.132 51.876 ;
        RECT 48.158 51.834 65.086 51.922 ;
        RECT 57.082 42.91 74.023 42.985 ;
        RECT 65.04 34.952 65.086 51.922 ;
        RECT 48.112 51.88 65.04 51.968 ;
        RECT 57.128 42.864 74.069 42.939 ;
        RECT 64.994 34.998 65.04 51.968 ;
        RECT 48.066 51.926 64.994 52.014 ;
        RECT 57.174 42.818 74.115 42.893 ;
        RECT 64.948 35.044 64.994 52.014 ;
        RECT 48.02 51.972 64.948 52.06 ;
        RECT 57.22 42.772 74.161 42.847 ;
        RECT 64.902 35.09 64.948 52.06 ;
        RECT 47.974 52.018 64.902 52.106 ;
        RECT 57.266 42.726 74.207 42.801 ;
        RECT 64.856 35.136 64.902 52.106 ;
        RECT 47.928 52.064 64.856 52.152 ;
        RECT 57.312 42.68 74.253 42.755 ;
        RECT 64.81 35.182 64.856 52.152 ;
        RECT 47.882 52.11 64.81 52.198 ;
        RECT 57.358 42.634 74.299 42.709 ;
        RECT 64.764 35.228 64.81 52.198 ;
        RECT 47.836 52.156 64.764 52.244 ;
        RECT 57.404 42.588 74.345 42.663 ;
        RECT 64.718 35.274 64.764 52.244 ;
        RECT 47.79 52.202 64.718 52.29 ;
        RECT 57.45 42.542 74.391 42.617 ;
        RECT 64.672 35.32 64.718 52.29 ;
        RECT 47.744 52.248 64.672 52.336 ;
        RECT 57.496 42.496 74.437 42.571 ;
        RECT 64.626 35.366 64.672 52.336 ;
        RECT 47.698 52.294 64.626 52.382 ;
        RECT 57.542 42.45 110 42.5 ;
        RECT 64.58 35.412 64.626 52.382 ;
        RECT 47.652 52.34 64.58 52.428 ;
        RECT 57.588 42.404 110 42.5 ;
        RECT 64.534 35.458 64.58 52.428 ;
        RECT 47.606 52.386 64.534 52.474 ;
        RECT 57.634 42.358 110 42.5 ;
        RECT 64.488 35.504 64.534 52.474 ;
        RECT 47.56 52.432 64.488 52.52 ;
        RECT 57.68 42.312 110 42.5 ;
        RECT 64.442 35.55 64.488 52.52 ;
        RECT 47.514 52.478 64.442 52.566 ;
        RECT 57.726 42.266 110 42.5 ;
        RECT 64.396 35.596 64.442 52.566 ;
        RECT 47.468 52.524 64.396 52.612 ;
        RECT 57.772 42.22 110 42.5 ;
        RECT 64.35 35.642 64.396 52.612 ;
        RECT 47.422 52.57 64.35 52.658 ;
        RECT 57.818 42.174 110 42.5 ;
        RECT 64.304 35.688 64.35 52.658 ;
        RECT 47.376 52.616 64.304 52.704 ;
        RECT 57.864 42.128 110 42.5 ;
        RECT 64.258 35.734 64.304 52.704 ;
        RECT 47.33 52.662 64.258 52.75 ;
        RECT 57.91 42.082 110 42.5 ;
        RECT 64.212 35.78 64.258 52.75 ;
        RECT 47.284 52.708 64.212 52.796 ;
        RECT 57.956 42.036 110 42.5 ;
        RECT 64.166 35.826 64.212 52.796 ;
        RECT 47.238 52.754 64.166 52.842 ;
        RECT 58.002 41.99 110 42.5 ;
        RECT 64.12 35.872 64.166 52.842 ;
        RECT 47.192 52.8 64.12 52.888 ;
        RECT 58.048 41.944 110 42.5 ;
        RECT 64.074 35.918 64.12 52.888 ;
        RECT 47.146 52.846 64.074 52.934 ;
        RECT 58.094 41.898 110 42.5 ;
        RECT 64.028 35.964 64.074 52.934 ;
        RECT 47.1 52.892 64.028 52.98 ;
        RECT 58.14 41.852 110 42.5 ;
        RECT 63.982 36.01 64.028 52.98 ;
        RECT 47.054 52.938 63.982 53.026 ;
        RECT 58.186 41.806 110 42.5 ;
        RECT 63.936 36.056 63.982 53.026 ;
        RECT 47.008 52.984 63.936 53.072 ;
        RECT 58.232 41.76 110 42.5 ;
        RECT 63.89 36.102 63.936 53.072 ;
        RECT 46.962 53.03 63.89 53.118 ;
        RECT 58.278 41.714 110 42.5 ;
        RECT 63.844 36.148 63.89 53.118 ;
        RECT 46.916 53.076 63.844 53.164 ;
        RECT 58.324 41.668 110 42.5 ;
        RECT 63.798 36.194 63.844 53.164 ;
        RECT 46.87 53.122 63.798 53.21 ;
        RECT 58.37 41.622 110 42.5 ;
        RECT 63.752 36.24 63.798 53.21 ;
        RECT 46.824 53.168 63.752 53.256 ;
        RECT 58.416 41.576 110 42.5 ;
        RECT 63.706 36.286 63.752 53.256 ;
        RECT 46.778 53.214 63.706 53.302 ;
        RECT 58.462 41.53 110 42.5 ;
        RECT 63.66 36.332 63.706 53.302 ;
        RECT 46.732 53.26 63.66 53.348 ;
        RECT 58.508 41.484 110 42.5 ;
        RECT 63.614 36.378 63.66 53.348 ;
        RECT 46.686 53.306 63.614 53.394 ;
        RECT 58.554 41.438 110 42.5 ;
        RECT 63.568 36.424 63.614 53.394 ;
        RECT 46.64 53.352 63.568 53.44 ;
        RECT 58.6 41.392 110 42.5 ;
        RECT 63.522 36.47 63.568 53.44 ;
        RECT 46.594 53.398 63.522 53.486 ;
        RECT 58.646 41.346 110 42.5 ;
        RECT 63.476 36.516 63.522 53.486 ;
        RECT 46.548 53.444 63.476 53.532 ;
        RECT 58.692 41.3 110 42.5 ;
        RECT 63.43 36.562 63.476 53.532 ;
        RECT 46.502 53.49 63.43 53.578 ;
        RECT 58.738 41.254 110 42.5 ;
        RECT 63.384 36.608 63.43 53.578 ;
        RECT 46.456 53.536 63.384 53.624 ;
        RECT 58.784 41.208 110 42.5 ;
        RECT 63.338 36.654 63.384 53.624 ;
        RECT 46.41 53.582 63.338 53.67 ;
        RECT 58.83 41.162 110 42.5 ;
        RECT 63.292 36.7 63.338 53.67 ;
        RECT 46.364 53.628 63.292 53.716 ;
        RECT 58.876 41.116 110 42.5 ;
        RECT 63.246 36.746 63.292 53.716 ;
        RECT 46.318 53.674 63.246 53.762 ;
        RECT 58.922 41.07 110 42.5 ;
        RECT 63.2 36.792 63.246 53.762 ;
        RECT 46.272 53.72 63.2 53.808 ;
        RECT 58.968 41.024 110 42.5 ;
        RECT 63.154 36.838 63.2 53.808 ;
        RECT 46.226 53.766 63.154 53.854 ;
        RECT 59.014 40.978 110 42.5 ;
        RECT 63.108 36.884 63.154 53.854 ;
        RECT 46.18 53.812 63.108 53.9 ;
        RECT 59.06 40.932 110 42.5 ;
        RECT 63.062 36.93 63.108 53.9 ;
        RECT 46.134 53.858 63.062 53.946 ;
        RECT 59.106 40.886 110 42.5 ;
        RECT 63.016 36.976 63.062 53.946 ;
        RECT 46.088 53.904 63.016 53.992 ;
        RECT 59.152 40.84 110 42.5 ;
        RECT 62.97 37.022 63.016 53.992 ;
        RECT 46.042 53.95 62.97 54.038 ;
        RECT 59.198 40.794 110 42.5 ;
        RECT 62.924 37.068 62.97 54.038 ;
        RECT 45.996 53.996 62.924 54.084 ;
        RECT 59.244 40.748 110 42.5 ;
        RECT 62.878 37.114 62.924 54.084 ;
        RECT 45.95 54.042 62.878 54.13 ;
        RECT 59.29 40.702 110 42.5 ;
        RECT 62.832 37.16 62.878 54.13 ;
        RECT 45.904 54.088 62.832 54.176 ;
        RECT 59.336 40.656 110 42.5 ;
        RECT 62.786 37.206 62.832 54.176 ;
        RECT 45.858 54.134 62.786 54.222 ;
        RECT 59.382 40.61 110 42.5 ;
        RECT 62.74 37.252 62.786 54.222 ;
        RECT 45.812 54.18 62.74 54.268 ;
        RECT 59.428 40.564 110 42.5 ;
        RECT 62.694 37.298 62.74 54.268 ;
        RECT 45.766 54.226 62.694 54.314 ;
        RECT 59.474 40.518 110 42.5 ;
        RECT 62.648 37.344 62.694 54.314 ;
        RECT 45.72 54.272 62.648 54.36 ;
        RECT 59.52 40.472 110 42.5 ;
        RECT 62.602 37.39 62.648 54.36 ;
        RECT 45.674 54.318 62.602 54.406 ;
        RECT 59.566 40.426 110 42.5 ;
        RECT 62.556 37.436 62.602 54.406 ;
        RECT 45.628 54.364 62.556 54.452 ;
        RECT 59.612 40.38 110 42.5 ;
        RECT 62.51 37.482 62.556 54.452 ;
        RECT 45.582 54.41 62.51 54.498 ;
        RECT 59.658 40.334 110 42.5 ;
        RECT 62.464 37.528 62.51 54.498 ;
        RECT 45.536 54.456 62.464 54.544 ;
        RECT 59.704 40.288 110 42.5 ;
        RECT 62.418 37.574 62.464 54.544 ;
        RECT 45.49 54.502 62.418 54.59 ;
        RECT 59.75 40.242 110 42.5 ;
        RECT 62.372 37.62 62.418 54.59 ;
        RECT 45.444 54.548 62.372 54.636 ;
        RECT 59.796 40.196 110 42.5 ;
        RECT 62.326 37.666 62.372 54.636 ;
        RECT 45.398 54.594 62.326 54.682 ;
        RECT 59.842 40.15 110 42.5 ;
        RECT 62.28 37.712 62.326 54.682 ;
        RECT 45.352 54.64 62.28 54.728 ;
        RECT 59.888 40.104 110 42.5 ;
        RECT 62.234 37.758 62.28 54.728 ;
        RECT 45.306 54.686 62.234 54.774 ;
        RECT 59.934 40.058 110 42.5 ;
        RECT 62.188 37.804 62.234 54.774 ;
        RECT 45.26 54.732 62.188 54.82 ;
        RECT 59.98 40.012 110 42.5 ;
        RECT 62.142 37.85 62.188 54.82 ;
        RECT 45.214 54.778 62.142 54.866 ;
        RECT 60.026 39.966 110 42.5 ;
        RECT 62.096 37.896 62.142 54.866 ;
        RECT 45.168 54.824 62.096 54.912 ;
        RECT 60.072 39.92 110 42.5 ;
        RECT 62.05 37.942 62.096 54.912 ;
        RECT 45.122 54.87 62.05 54.958 ;
        RECT 60.118 39.874 110 42.5 ;
        RECT 62.004 37.988 62.05 54.958 ;
        RECT 45.076 54.916 62.004 55.004 ;
        RECT 60.164 39.828 110 42.5 ;
        RECT 61.958 38.034 62.004 55.004 ;
        RECT 45.03 54.962 61.958 55.05 ;
        RECT 60.21 39.782 110 42.5 ;
        RECT 61.912 38.08 61.958 55.05 ;
        RECT 44.984 55.008 61.912 55.096 ;
        RECT 60.256 39.736 110 42.5 ;
        RECT 61.866 38.126 61.912 55.096 ;
        RECT 44.938 55.054 61.866 55.142 ;
        RECT 60.302 39.69 110 42.5 ;
        RECT 61.82 38.172 61.866 55.142 ;
        RECT 44.892 55.1 61.82 55.188 ;
        RECT 60.348 39.644 110 42.5 ;
        RECT 61.774 38.218 61.82 55.188 ;
        RECT 44.846 55.146 61.774 55.234 ;
        RECT 60.394 39.598 110 42.5 ;
        RECT 61.728 38.264 61.774 55.234 ;
        RECT 44.8 55.192 61.728 55.28 ;
        RECT 60.44 39.552 110 42.5 ;
        RECT 61.682 38.31 61.728 55.28 ;
        RECT 44.754 55.238 61.682 55.326 ;
        RECT 60.486 39.506 110 42.5 ;
        RECT 61.636 38.356 61.682 55.326 ;
        RECT 44.708 55.284 61.636 55.372 ;
        RECT 60.532 39.46 110 42.5 ;
        RECT 61.59 38.402 61.636 55.372 ;
        RECT 44.662 55.33 61.59 55.418 ;
        RECT 60.578 39.414 110 42.5 ;
        RECT 61.544 38.448 61.59 55.418 ;
        RECT 44.616 55.376 61.544 55.464 ;
        RECT 60.624 39.368 110 42.5 ;
        RECT 61.498 38.494 61.544 55.464 ;
        RECT 44.57 55.422 61.498 55.51 ;
        RECT 60.67 39.322 110 42.5 ;
        RECT 61.452 38.54 61.498 55.51 ;
        RECT 44.524 55.468 61.452 55.556 ;
        RECT 60.716 39.276 110 42.5 ;
        RECT 61.406 38.586 61.452 55.556 ;
        RECT 44.478 55.514 61.406 55.602 ;
        RECT 60.762 39.23 110 42.5 ;
        RECT 61.36 38.632 61.406 55.602 ;
        RECT 44.432 55.56 61.36 55.648 ;
        RECT 60.808 39.184 110 42.5 ;
        RECT 61.314 38.678 61.36 55.648 ;
        RECT 44.386 55.606 61.314 55.694 ;
        RECT 60.854 39.138 110 42.5 ;
        RECT 61.268 38.724 61.314 55.694 ;
        RECT 44.34 55.652 61.268 55.74 ;
        RECT 60.9 39.092 110 42.5 ;
        RECT 61.222 38.77 61.268 55.74 ;
        RECT 44.294 55.698 61.222 55.786 ;
        RECT 60.946 39.046 110 42.5 ;
        RECT 61.176 38.816 61.222 55.786 ;
        RECT 44.248 55.744 61.176 55.832 ;
        RECT 60.992 39 110 42.5 ;
        RECT 61.13 38.862 61.176 55.832 ;
        RECT 44.202 55.79 61.13 55.878 ;
        RECT 61.038 38.954 110 42.5 ;
        RECT 61.084 38.908 61.13 55.878 ;
        RECT 44.156 55.836 61.084 55.924 ;
        RECT 44.11 55.882 61.038 55.97 ;
        RECT 44.064 55.928 60.992 56.016 ;
        RECT 44.018 55.974 60.946 56.062 ;
        RECT 43.972 56.02 60.9 56.108 ;
        RECT 43.926 56.066 60.854 56.154 ;
        RECT 43.88 56.112 60.808 56.2 ;
        RECT 43.834 56.158 60.762 56.246 ;
        RECT 43.788 56.204 60.716 56.292 ;
        RECT 43.742 56.25 60.67 56.338 ;
        RECT 43.696 56.296 60.624 56.384 ;
        RECT 43.65 56.342 60.578 56.43 ;
        RECT 43.604 56.388 60.532 56.476 ;
        RECT 43.558 56.434 60.486 56.522 ;
        RECT 43.512 56.48 60.44 56.568 ;
        RECT 43.466 56.526 60.394 56.614 ;
        RECT 43.42 56.572 60.348 56.66 ;
        RECT 43.374 56.618 60.302 56.706 ;
        RECT 43.328 56.664 60.256 56.752 ;
        RECT 43.282 56.71 60.21 56.798 ;
        RECT 43.236 56.756 60.164 56.844 ;
        RECT 43.19 56.802 60.118 56.89 ;
        RECT 43.144 56.848 60.072 56.936 ;
        RECT 43.098 56.894 60.026 56.982 ;
        RECT 43.052 56.94 59.98 57.028 ;
        RECT 43.006 56.986 59.934 57.074 ;
        RECT 42.96 57.032 59.888 57.12 ;
        RECT 42.914 57.078 59.842 57.166 ;
        RECT 42.868 57.124 59.796 57.212 ;
        RECT 42.822 57.17 59.75 57.258 ;
        RECT 42.776 57.216 59.704 57.304 ;
        RECT 42.73 57.262 59.658 57.35 ;
        RECT 42.684 57.308 59.612 57.396 ;
        RECT 42.638 57.354 59.566 57.442 ;
        RECT 42.592 57.4 59.52 57.488 ;
        RECT 42.5 57.492 59.474 57.534 ;
        RECT 42.546 57.446 59.474 57.534 ;
        RECT 42.46 57.535 59.428 57.58 ;
        RECT 42.414 57.578 59.382 57.626 ;
        RECT 42.368 57.624 59.336 57.672 ;
        RECT 42.322 57.67 59.29 57.718 ;
        RECT 42.276 57.716 59.244 57.764 ;
        RECT 42.23 57.762 59.198 57.81 ;
        RECT 42.184 57.808 59.152 57.856 ;
        RECT 42.138 57.854 59.106 57.902 ;
        RECT 42.092 57.9 59.06 57.948 ;
        RECT 42.046 57.946 59.014 57.994 ;
        RECT 42 57.992 58.968 58.04 ;
        RECT 41.954 58.038 58.922 58.086 ;
        RECT 41.908 58.084 58.876 58.132 ;
        RECT 41.862 58.13 58.83 58.178 ;
        RECT 41.816 58.176 58.784 58.224 ;
        RECT 41.77 58.222 58.738 58.27 ;
        RECT 41.724 58.268 58.692 58.316 ;
        RECT 41.678 58.314 58.646 58.362 ;
        RECT 41.632 58.36 58.6 58.408 ;
        RECT 41.586 58.406 58.554 58.454 ;
        RECT 41.54 58.452 58.508 58.5 ;
        RECT 41.494 58.498 58.462 58.546 ;
        RECT 41.448 58.544 58.416 58.592 ;
        RECT 41.402 58.59 58.37 58.638 ;
        RECT 41.356 58.636 58.324 58.684 ;
        RECT 41.31 58.682 58.278 58.73 ;
        RECT 41.264 58.728 58.232 58.776 ;
        RECT 41.218 58.774 58.186 58.822 ;
        RECT 41.172 58.82 58.14 58.868 ;
        RECT 41.126 58.866 58.094 58.914 ;
        RECT 41.08 58.912 58.048 58.96 ;
        RECT 41.034 58.958 58.002 59.006 ;
        RECT 40.988 59.004 57.956 59.052 ;
        RECT 40.942 59.05 57.91 59.098 ;
        RECT 40.896 59.096 57.864 59.144 ;
        RECT 40.85 59.142 57.818 59.19 ;
        RECT 40.804 59.188 57.772 59.236 ;
        RECT 40.758 59.234 57.726 59.282 ;
        RECT 40.712 59.28 57.68 59.328 ;
        RECT 40.666 59.326 57.634 59.374 ;
        RECT 40.62 59.372 57.588 59.42 ;
        RECT 40.574 59.418 57.542 59.466 ;
        RECT 40.528 59.464 57.496 59.512 ;
        RECT 40.482 59.51 57.45 59.558 ;
        RECT 40.436 59.556 57.404 59.604 ;
        RECT 40.39 59.602 57.358 59.65 ;
        RECT 40.344 59.648 57.312 59.696 ;
        RECT 40.298 59.694 57.266 59.742 ;
        RECT 40.252 59.74 57.22 59.788 ;
        RECT 40.206 59.786 57.174 59.834 ;
        RECT 40.16 59.832 57.128 59.88 ;
        RECT 40.114 59.878 57.082 59.926 ;
        RECT 40.068 59.924 57.036 59.972 ;
        RECT 40.022 59.97 56.99 60.018 ;
        RECT 39.976 60.016 56.944 60.064 ;
        RECT 39.93 60.062 56.898 60.11 ;
        RECT 39.884 60.108 56.852 60.156 ;
        RECT 39.838 60.154 56.806 60.202 ;
        RECT 39.792 60.2 56.76 60.248 ;
        RECT 39.746 60.246 56.714 60.294 ;
        RECT 39.7 60.292 56.668 60.34 ;
        RECT 39.654 60.338 56.622 60.386 ;
        RECT 39.608 60.384 56.576 60.432 ;
        RECT 39.562 60.43 56.53 60.478 ;
        RECT 39.516 60.476 56.484 60.524 ;
        RECT 39.47 60.522 56.438 60.57 ;
        RECT 39.424 60.568 56.392 60.616 ;
        RECT 39.378 60.614 56.346 60.662 ;
        RECT 39.332 60.66 56.3 60.708 ;
        RECT 39.286 60.706 56.254 60.754 ;
        RECT 39.24 60.752 56.208 60.8 ;
        RECT 39.194 60.798 56.162 60.846 ;
        RECT 39.148 60.844 56.116 60.892 ;
        RECT 39.102 60.89 56.07 60.938 ;
        RECT 39.056 60.936 56.024 60.984 ;
        RECT 39.01 60.982 55.978 61.03 ;
        RECT 38.964 61.028 55.932 61.076 ;
        RECT 38.918 61.074 55.886 61.122 ;
        RECT 38.872 61.12 55.84 61.168 ;
        RECT 38.826 61.166 55.794 61.214 ;
        RECT 38.78 61.212 55.748 61.26 ;
        RECT 38.734 61.258 55.702 61.306 ;
        RECT 38.688 61.304 55.656 61.352 ;
        RECT 38.642 61.35 55.61 61.398 ;
        RECT 38.596 61.396 55.564 61.444 ;
        RECT 38.55 61.442 55.518 61.49 ;
        RECT 38.504 61.488 55.472 61.536 ;
        RECT 38.458 61.534 55.426 61.582 ;
        RECT 38.412 61.58 55.38 61.628 ;
        RECT 38.366 61.626 55.334 61.674 ;
        RECT 38.32 61.672 55.288 61.72 ;
        RECT 38.274 61.718 55.242 61.766 ;
        RECT 38.228 61.764 55.196 61.812 ;
        RECT 38.182 61.81 55.15 61.858 ;
        RECT 38.136 61.856 55.104 61.904 ;
        RECT 38.09 61.902 55.058 61.95 ;
        RECT 38.044 61.948 55.012 61.996 ;
        RECT 37.998 61.994 54.966 62.042 ;
        RECT 37.952 62.04 54.92 62.088 ;
        RECT 37.906 62.086 54.874 62.134 ;
        RECT 37.86 62.132 54.828 62.18 ;
        RECT 37.814 62.178 54.782 62.226 ;
        RECT 37.768 62.224 54.736 62.272 ;
        RECT 37.722 62.27 54.69 62.318 ;
        RECT 37.676 62.316 54.644 62.364 ;
        RECT 37.63 62.362 54.598 62.41 ;
        RECT 37.584 62.408 54.552 62.456 ;
        RECT 37.538 62.454 54.506 62.502 ;
        RECT 37.492 62.5 54.46 62.548 ;
        RECT 37.446 62.546 54.414 62.594 ;
        RECT 37.4 62.592 54.368 62.64 ;
        RECT 37.354 62.638 54.322 62.686 ;
        RECT 37.308 62.684 54.276 62.732 ;
        RECT 37.262 62.73 54.23 62.778 ;
        RECT 37.216 62.776 54.184 62.824 ;
        RECT 37.17 62.822 54.138 62.87 ;
        RECT 37.124 62.868 54.092 62.916 ;
        RECT 37.078 62.914 54.046 62.962 ;
        RECT 37.032 62.96 54 63.008 ;
        RECT 36.986 63.006 53.954 63.054 ;
        RECT 36.94 63.052 53.908 63.1 ;
        RECT 36.894 63.098 53.862 63.146 ;
        RECT 36.848 63.144 53.816 63.192 ;
        RECT 36.802 63.19 53.77 63.238 ;
        RECT 36.756 63.236 53.724 63.284 ;
        RECT 36.71 63.282 53.678 63.33 ;
        RECT 36.664 63.328 53.632 63.376 ;
        RECT 36.618 63.374 53.586 63.422 ;
        RECT 36.572 63.42 53.54 63.468 ;
        RECT 36.526 63.466 53.494 63.514 ;
        RECT 36.48 63.512 53.448 63.56 ;
        RECT 36.434 63.558 53.402 63.606 ;
        RECT 36.388 63.604 53.356 63.652 ;
        RECT 36.342 63.65 53.31 63.698 ;
        RECT 36.296 63.696 53.264 63.744 ;
        RECT 36.25 63.742 53.218 63.79 ;
        RECT 36.204 63.788 53.172 63.836 ;
        RECT 36.158 63.834 53.126 63.882 ;
        RECT 36.112 63.88 53.08 63.928 ;
        RECT 36.066 63.926 53.034 63.974 ;
        RECT 36.02 63.972 52.988 64.02 ;
        RECT 35.974 64.018 52.942 64.066 ;
        RECT 35.928 64.064 52.896 64.112 ;
        RECT 35.882 64.11 52.85 64.158 ;
        RECT 35.836 64.156 52.804 64.204 ;
        RECT 35.79 64.202 52.758 64.25 ;
        RECT 35.744 64.248 52.712 64.296 ;
        RECT 35.698 64.294 52.666 64.342 ;
        RECT 35.652 64.34 52.62 64.388 ;
        RECT 35.606 64.386 52.574 64.434 ;
        RECT 35.56 64.432 52.528 64.48 ;
        RECT 35.514 64.478 52.482 64.526 ;
        RECT 35.468 64.524 52.436 64.572 ;
        RECT 35.422 64.57 52.39 64.618 ;
        RECT 35.376 64.616 52.344 64.664 ;
        RECT 35.33 64.662 52.298 64.71 ;
        RECT 35.284 64.708 52.252 64.756 ;
        RECT 35.238 64.754 52.206 64.802 ;
        RECT 35.192 64.8 52.16 64.848 ;
        RECT 35.146 64.846 52.114 64.894 ;
        RECT 35.1 64.892 52.068 64.94 ;
        RECT 35.054 64.938 52.022 64.986 ;
        RECT 35.008 64.984 51.976 65.032 ;
        RECT 34.962 65.03 51.93 65.078 ;
        RECT 34.916 65.076 51.884 65.124 ;
        RECT 34.87 65.122 51.838 65.17 ;
        RECT 34.824 65.168 51.792 65.216 ;
        RECT 34.778 65.214 51.746 65.262 ;
        RECT 34.732 65.26 51.7 65.308 ;
        RECT 34.686 65.306 51.654 65.354 ;
        RECT 34.64 65.352 51.608 65.4 ;
        RECT 34.594 65.398 51.562 65.446 ;
        RECT 34.548 65.444 51.516 65.492 ;
        RECT 34.502 65.49 51.47 65.538 ;
        RECT 34.456 65.536 51.424 65.584 ;
        RECT 34.41 65.582 51.378 65.63 ;
        RECT 34.364 65.628 51.332 65.676 ;
        RECT 34.318 65.674 51.286 65.722 ;
        RECT 34.272 65.72 51.24 65.768 ;
        RECT 34.226 65.766 51.194 65.814 ;
        RECT 34.18 65.812 51.148 65.86 ;
        RECT 34.134 65.858 51.102 65.906 ;
        RECT 34.088 65.904 51.056 65.952 ;
        RECT 34.042 65.95 51.01 65.998 ;
        RECT 33.996 65.996 50.964 66.044 ;
        RECT 33.95 66.042 50.918 66.09 ;
        RECT 33.904 66.088 50.872 66.136 ;
        RECT 33.858 66.134 50.826 66.182 ;
        RECT 33.812 66.18 50.78 66.228 ;
        RECT 33.766 66.226 50.734 66.274 ;
        RECT 33.72 66.272 50.688 66.32 ;
        RECT 33.674 66.318 50.642 66.366 ;
        RECT 33.628 66.364 50.596 66.412 ;
        RECT 33.582 66.41 50.55 66.458 ;
        RECT 33.536 66.456 50.504 66.504 ;
        RECT 33.49 66.502 50.458 66.55 ;
        RECT 33.444 66.548 50.412 66.596 ;
        RECT 33.398 66.594 50.366 66.642 ;
        RECT 33.352 66.64 50.32 66.688 ;
        RECT 33.306 66.686 50.274 66.734 ;
        RECT 33.26 66.732 50.228 66.78 ;
        RECT 33.214 66.778 50.182 66.826 ;
        RECT 33.168 66.824 50.136 66.872 ;
        RECT 33.122 66.87 50.09 66.918 ;
        RECT 33.076 66.916 50.044 66.964 ;
        RECT 33.03 66.962 49.998 67.01 ;
        RECT 32.984 67.008 49.952 67.056 ;
        RECT 32.938 67.054 49.906 67.102 ;
        RECT 32.892 67.1 49.86 67.148 ;
        RECT 32.846 67.146 49.814 67.194 ;
        RECT 32.8 67.192 49.768 67.24 ;
        RECT 32.754 67.238 49.722 67.286 ;
        RECT 32.708 67.284 49.676 67.332 ;
        RECT 32.662 67.33 49.63 67.378 ;
        RECT 32.616 67.376 49.584 67.424 ;
        RECT 32.57 67.422 49.538 67.47 ;
        RECT 32.524 67.468 49.492 67.516 ;
        RECT 32.478 67.514 49.446 67.562 ;
        RECT 32.432 67.56 49.4 67.608 ;
        RECT 32.386 67.606 49.354 67.654 ;
        RECT 32.34 67.652 49.308 67.7 ;
        RECT 32.294 67.698 49.262 67.746 ;
        RECT 32.248 67.744 49.216 67.792 ;
        RECT 32.202 67.79 49.17 67.838 ;
        RECT 32.156 67.836 49.124 67.884 ;
        RECT 32.11 67.882 49.078 67.93 ;
        RECT 32.064 67.928 49.032 67.976 ;
        RECT 32.018 67.974 48.986 68.022 ;
        RECT 31.972 68.02 48.94 68.068 ;
        RECT 31.926 68.066 48.894 68.114 ;
        RECT 31.88 68.112 48.848 68.16 ;
        RECT 31.834 68.158 48.802 68.206 ;
        RECT 31.788 68.204 48.756 68.252 ;
        RECT 31.742 68.25 48.71 68.298 ;
        RECT 31.696 68.296 48.664 68.344 ;
        RECT 31.65 68.342 48.618 68.39 ;
        RECT 31.604 68.388 48.572 68.436 ;
        RECT 31.558 68.434 48.526 68.482 ;
        RECT 31.512 68.48 48.48 68.528 ;
        RECT 31.466 68.526 48.434 68.574 ;
        RECT 31.42 68.572 48.388 68.62 ;
        RECT 31.374 68.618 48.342 68.666 ;
        RECT 31.328 68.664 48.296 68.712 ;
        RECT 31.282 68.71 48.25 68.758 ;
        RECT 31.236 68.756 48.204 68.804 ;
        RECT 31.19 68.802 48.158 68.85 ;
        RECT 31.144 68.848 48.112 68.896 ;
        RECT 31.098 68.894 48.066 68.942 ;
        RECT 31.052 68.94 48.02 68.988 ;
        RECT 31.006 68.986 47.974 69.034 ;
        RECT 30.96 69.032 47.928 69.08 ;
        RECT 30.914 69.078 47.882 69.126 ;
        RECT 30.868 69.124 47.836 69.172 ;
        RECT 30.822 69.17 47.79 69.218 ;
        RECT 30.776 69.216 47.744 69.264 ;
        RECT 30.73 69.262 47.698 69.31 ;
        RECT 30.684 69.308 47.652 69.356 ;
        RECT 30.638 69.354 47.606 69.402 ;
        RECT 30.592 69.4 47.56 69.448 ;
        RECT 30.546 69.446 47.514 69.494 ;
        RECT 30.5 69.492 47.468 69.54 ;
        RECT 30.5 69.492 47.422 69.586 ;
        RECT 30.5 69.492 47.376 69.632 ;
        RECT 30.5 69.492 47.33 69.678 ;
        RECT 30.5 69.492 47.284 69.724 ;
        RECT 30.5 69.492 47.238 69.77 ;
        RECT 30.5 69.492 47.192 69.816 ;
        RECT 30.5 69.492 47.146 69.862 ;
        RECT 30.5 69.492 47.1 69.908 ;
        RECT 30.5 69.492 47.054 69.954 ;
        RECT 30.5 69.492 47.008 70 ;
        RECT 30.5 69.492 46.962 70.046 ;
        RECT 30.5 69.492 46.916 70.092 ;
        RECT 30.5 69.492 46.87 70.138 ;
        RECT 30.5 69.492 46.824 70.184 ;
        RECT 30.5 69.492 46.778 70.23 ;
        RECT 30.5 69.492 46.732 70.276 ;
        RECT 30.5 69.492 46.686 70.322 ;
        RECT 30.5 69.492 46.64 70.368 ;
        RECT 30.5 69.492 46.594 70.414 ;
        RECT 30.5 69.492 46.548 70.46 ;
        RECT 30.5 69.492 46.502 70.506 ;
        RECT 30.5 69.492 46.456 70.552 ;
        RECT 30.5 69.492 46.41 70.598 ;
        RECT 30.5 69.492 46.364 70.644 ;
        RECT 30.5 69.492 46.318 70.69 ;
        RECT 30.5 69.492 46.272 70.736 ;
        RECT 30.5 69.492 46.226 70.782 ;
        RECT 30.5 69.492 46.18 70.828 ;
        RECT 30.5 69.492 46.134 70.874 ;
        RECT 30.5 69.492 46.088 70.92 ;
        RECT 30.5 69.492 46.042 70.966 ;
        RECT 30.5 69.492 45.996 71.012 ;
        RECT 30.5 69.492 45.95 71.058 ;
        RECT 30.5 69.492 45.904 71.104 ;
        RECT 30.5 69.492 45.858 71.15 ;
        RECT 30.5 69.492 45.812 71.196 ;
        RECT 30.5 69.492 45.766 71.242 ;
        RECT 30.5 69.492 45.72 71.288 ;
        RECT 30.5 69.492 45.674 71.334 ;
        RECT 30.5 69.492 45.628 71.38 ;
        RECT 30.5 69.492 45.582 71.426 ;
        RECT 30.5 69.492 45.536 71.472 ;
        RECT 30.5 69.492 45.49 71.518 ;
        RECT 30.5 69.492 45.444 71.564 ;
        RECT 30.5 69.492 45.398 71.61 ;
        RECT 30.5 69.492 45.352 71.656 ;
        RECT 30.5 69.492 45.306 71.702 ;
        RECT 30.5 69.492 45.26 71.748 ;
        RECT 30.5 69.492 45.214 71.794 ;
        RECT 30.5 69.492 45.168 71.84 ;
        RECT 30.5 69.492 45.122 71.886 ;
        RECT 30.5 69.492 45.076 71.932 ;
        RECT 30.5 69.492 45.03 71.978 ;
        RECT 30.5 69.492 44.984 72.024 ;
        RECT 30.5 69.492 44.938 72.07 ;
        RECT 30.5 69.492 44.892 72.116 ;
        RECT 30.5 69.492 44.846 72.162 ;
        RECT 30.5 69.492 44.8 72.208 ;
        RECT 30.5 69.492 44.754 72.254 ;
        RECT 30.5 69.492 44.708 72.3 ;
        RECT 30.5 69.492 44.662 72.346 ;
        RECT 30.5 69.492 44.616 72.392 ;
        RECT 30.5 69.492 44.57 72.438 ;
        RECT 30.5 69.492 44.524 72.484 ;
        RECT 30.5 69.492 44.478 72.53 ;
        RECT 30.5 69.492 44.432 72.576 ;
        RECT 30.5 69.492 44.386 72.622 ;
        RECT 30.5 69.492 44.34 72.668 ;
        RECT 30.5 69.492 44.294 72.714 ;
        RECT 30.5 69.492 44.248 72.76 ;
        RECT 30.5 69.492 44.202 72.806 ;
        RECT 30.5 69.492 44.156 72.852 ;
        RECT 30.5 69.492 44.11 72.898 ;
        RECT 30.5 69.492 44.064 72.944 ;
        RECT 30.5 69.492 44.018 72.99 ;
        RECT 30.5 69.492 43.972 73.036 ;
        RECT 30.5 69.492 43.926 73.082 ;
        RECT 30.5 69.492 43.88 73.128 ;
        RECT 30.5 69.492 43.834 73.174 ;
        RECT 30.5 69.492 43.788 73.22 ;
        RECT 30.5 69.492 43.742 73.266 ;
        RECT 30.5 69.492 43.696 73.312 ;
        RECT 30.5 69.492 43.65 73.358 ;
        RECT 30.5 69.492 43.604 73.404 ;
        RECT 30.5 69.492 43.558 73.45 ;
        RECT 30.5 69.492 43.512 73.496 ;
        RECT 30.5 69.492 43.466 73.542 ;
        RECT 30.5 69.492 43.42 73.588 ;
        RECT 30.5 69.492 43.374 73.634 ;
        RECT 30.5 69.492 43.328 73.68 ;
        RECT 30.5 69.492 43.282 73.726 ;
        RECT 30.5 69.492 43.236 73.772 ;
        RECT 30.5 69.492 43.19 73.818 ;
        RECT 30.5 69.492 43.144 73.864 ;
        RECT 30.5 69.492 43.098 73.91 ;
        RECT 30.5 69.492 43.052 73.956 ;
        RECT 30.5 69.492 43.006 74.002 ;
        RECT 30.5 69.492 42.96 74.048 ;
        RECT 30.5 69.492 42.914 74.094 ;
        RECT 30.5 69.492 42.868 74.14 ;
        RECT 30.5 69.492 42.822 74.186 ;
        RECT 30.5 69.492 42.776 74.232 ;
        RECT 30.5 69.492 42.73 74.278 ;
        RECT 30.5 69.492 42.684 74.324 ;
        RECT 30.5 69.492 42.638 74.37 ;
        RECT 30.5 69.492 42.592 74.416 ;
        RECT 30.5 69.492 42.546 74.462 ;
        RECT 30.5 69.492 42.5 110 ;
        RECT 76.265 44 110 56 ;
        RECT 59.312 60.93 76.265 60.983 ;
        RECT 59.358 60.884 76.311 60.947 ;
        RECT 76.24 44.012 76.265 60.983 ;
        RECT 59.404 60.838 76.357 60.901 ;
        RECT 76.194 44.048 76.24 61.018 ;
        RECT 59.266 60.976 76.194 61.064 ;
        RECT 59.45 60.792 76.403 60.855 ;
        RECT 76.148 44.094 76.194 61.064 ;
        RECT 59.22 61.022 76.148 61.11 ;
        RECT 59.496 60.746 76.449 60.809 ;
        RECT 76.102 44.14 76.148 61.11 ;
        RECT 59.174 61.068 76.102 61.156 ;
        RECT 59.542 60.7 76.495 60.763 ;
        RECT 76.056 44.186 76.102 61.156 ;
        RECT 59.128 61.114 76.056 61.202 ;
        RECT 59.588 60.654 76.541 60.717 ;
        RECT 76.01 44.232 76.056 61.202 ;
        RECT 59.082 61.16 76.01 61.248 ;
        RECT 59.634 60.608 76.587 60.671 ;
        RECT 75.964 44.278 76.01 61.248 ;
        RECT 59.036 61.206 75.964 61.294 ;
        RECT 59.68 60.562 76.633 60.625 ;
        RECT 75.918 44.324 75.964 61.294 ;
        RECT 58.99 61.252 75.918 61.34 ;
        RECT 59.726 60.516 76.679 60.579 ;
        RECT 75.872 44.37 75.918 61.34 ;
        RECT 58.944 61.298 75.872 61.386 ;
        RECT 59.772 60.47 76.725 60.533 ;
        RECT 75.826 44.416 75.872 61.386 ;
        RECT 58.898 61.344 75.826 61.432 ;
        RECT 59.818 60.424 76.771 60.487 ;
        RECT 75.78 44.462 75.826 61.432 ;
        RECT 58.852 61.39 75.78 61.478 ;
        RECT 59.864 60.378 76.817 60.441 ;
        RECT 75.734 44.508 75.78 61.478 ;
        RECT 58.806 61.436 75.734 61.524 ;
        RECT 59.91 60.332 76.863 60.395 ;
        RECT 75.688 44.554 75.734 61.524 ;
        RECT 58.76 61.482 75.688 61.57 ;
        RECT 59.956 60.286 76.909 60.349 ;
    END
  END VDDIO
  PIN VSS
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8e-05 LAYER MET4 ;
    ANTENNAPARTIALMETALAREA 4.8e-05 LAYER MET3 ;
    ANTENNAPARTIALMETALAREA 4.8e-05 LAYER MET5 ;
    ANTENNAPARTIALMETALAREA 4.8e-05 LAYER MET2 ;
    ANTENNAPARTIALCUTAREA 1.5876 LAYER VIA4 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 2.3328 LAYER VIA2 ;
    PORT
      LAYER MET5 ;
        RECT 99.55 91 110 98 ;
        RECT 91 99.527 100.884 99.589 ;
        RECT 91 99.527 100.838 99.635 ;
        RECT 91 99.527 100.792 99.681 ;
        RECT 91 99.527 100.746 99.727 ;
        RECT 91 99.527 100.7 99.773 ;
        RECT 91 99.527 100.654 99.819 ;
        RECT 91 99.527 100.608 99.865 ;
        RECT 91 99.527 100.562 99.911 ;
        RECT 91 99.527 100.516 99.957 ;
        RECT 91 99.527 100.47 100.003 ;
        RECT 91 99.527 100.424 100.049 ;
        RECT 91 99.527 100.378 100.095 ;
        RECT 91 99.527 100.332 100.141 ;
        RECT 91 99.527 100.286 100.187 ;
        RECT 91 99.527 100.24 100.233 ;
        RECT 91 99.527 100.194 100.279 ;
        RECT 91 99.527 100.148 100.325 ;
        RECT 91 99.527 100.102 100.371 ;
        RECT 91 99.527 100.056 100.417 ;
        RECT 91 99.527 100.01 100.463 ;
        RECT 91 99.527 99.964 100.509 ;
        RECT 91 99.527 99.918 100.555 ;
        RECT 91 99.527 99.872 100.601 ;
        RECT 91 99.527 99.826 100.647 ;
        RECT 91 99.527 99.78 100.693 ;
        RECT 91 99.527 99.734 100.739 ;
        RECT 91 99.527 99.688 100.785 ;
        RECT 91 99.527 99.642 100.831 ;
        RECT 91 99.527 99.596 100.877 ;
        RECT 91.046 99.481 100.93 99.543 ;
        RECT 99.518 91.016 99.55 100.916 ;
        RECT 91.092 99.435 100.976 99.497 ;
        RECT 99.472 91.055 99.518 100.955 ;
        RECT 91.138 99.389 101.022 99.451 ;
        RECT 99.426 91.101 99.472 101.001 ;
        RECT 91.184 99.343 101.068 99.405 ;
        RECT 99.38 91.147 99.426 101.047 ;
        RECT 91.23 99.297 101.114 99.359 ;
        RECT 99.334 91.193 99.38 101.093 ;
        RECT 91.276 99.251 101.16 99.313 ;
        RECT 99.288 91.239 99.334 101.139 ;
        RECT 91.322 99.205 101.206 99.267 ;
        RECT 99.242 91.285 99.288 101.185 ;
        RECT 91.368 99.159 101.252 99.221 ;
        RECT 99.196 91.331 99.242 101.231 ;
        RECT 91.414 99.113 101.298 99.175 ;
        RECT 99.15 91.377 99.196 101.277 ;
        RECT 91.46 99.067 101.344 99.129 ;
        RECT 99.104 91.423 99.15 101.323 ;
        RECT 91.506 99.021 101.39 99.083 ;
        RECT 99.058 91.469 99.104 101.369 ;
        RECT 91.552 98.975 101.436 99.037 ;
        RECT 99.012 91.515 99.058 101.415 ;
        RECT 91.598 98.929 101.482 98.991 ;
        RECT 98.966 91.561 99.012 101.461 ;
        RECT 91.644 98.883 101.528 98.945 ;
        RECT 98.92 91.607 98.966 101.507 ;
        RECT 91.69 98.837 101.574 98.899 ;
        RECT 98.874 91.653 98.92 101.553 ;
        RECT 91.736 98.791 101.62 98.853 ;
        RECT 98.828 91.699 98.874 101.599 ;
        RECT 91.782 98.745 101.666 98.807 ;
        RECT 98.782 91.745 98.828 101.645 ;
        RECT 91.828 98.699 101.712 98.761 ;
        RECT 98.736 91.791 98.782 101.691 ;
        RECT 91.874 98.653 101.758 98.715 ;
        RECT 98.69 91.837 98.736 101.737 ;
        RECT 91.92 98.607 101.804 98.669 ;
        RECT 98.644 91.883 98.69 101.783 ;
        RECT 91.966 98.561 101.85 98.623 ;
        RECT 98.598 91.929 98.644 101.829 ;
        RECT 92.012 98.515 101.896 98.577 ;
        RECT 98.552 91.975 98.598 101.875 ;
        RECT 92.058 98.469 101.942 98.531 ;
        RECT 98.506 92.021 98.552 101.921 ;
        RECT 92.104 98.423 101.988 98.485 ;
        RECT 98.46 92.067 98.506 101.967 ;
        RECT 92.15 98.377 102.034 98.439 ;
        RECT 98.414 92.113 98.46 102.013 ;
        RECT 92.196 98.331 102.08 98.393 ;
        RECT 98.368 92.159 98.414 102.059 ;
        RECT 92.242 98.285 102.126 98.347 ;
        RECT 98.322 92.205 98.368 102.105 ;
        RECT 92.288 98.239 102.172 98.301 ;
        RECT 98.276 92.251 98.322 102.151 ;
        RECT 92.334 98.193 102.218 98.255 ;
        RECT 98.23 92.297 98.276 102.197 ;
        RECT 92.38 98.147 102.264 98.209 ;
        RECT 98.184 92.343 98.23 102.243 ;
        RECT 92.426 98.101 102.31 98.163 ;
        RECT 98.138 92.389 98.184 102.289 ;
        RECT 92.472 98.055 102.356 98.117 ;
        RECT 98.092 92.435 98.138 102.335 ;
        RECT 92.518 98.009 102.402 98.071 ;
        RECT 98.046 92.481 98.092 102.381 ;
        RECT 92.564 97.963 102.448 98.024 ;
        RECT 98 92.527 98.046 102.427 ;
        RECT 91 99.527 98 110 ;
        RECT 92.61 97.917 110 98 ;
        RECT 97.992 92.554 98 110 ;
        RECT 92.656 97.871 110 98 ;
        RECT 97.946 92.581 98 110 ;
        RECT 92.702 97.825 110 98 ;
        RECT 97.9 92.627 98 110 ;
        RECT 92.748 97.779 110 98 ;
        RECT 97.854 92.673 98 110 ;
        RECT 92.794 97.733 110 98 ;
        RECT 97.808 92.719 98 110 ;
        RECT 92.84 97.687 110 98 ;
        RECT 97.762 92.765 98 110 ;
        RECT 92.886 97.641 110 98 ;
        RECT 97.716 92.811 98 110 ;
        RECT 92.932 97.595 110 98 ;
        RECT 97.67 92.857 98 110 ;
        RECT 92.978 97.549 110 98 ;
        RECT 97.624 92.903 98 110 ;
        RECT 93.024 97.503 110 98 ;
        RECT 97.578 92.949 98 110 ;
        RECT 93.07 97.457 110 98 ;
        RECT 97.532 92.995 98 110 ;
        RECT 93.116 97.411 110 98 ;
        RECT 97.486 93.041 98 110 ;
        RECT 93.162 97.365 110 98 ;
        RECT 97.44 93.087 98 110 ;
        RECT 93.208 97.319 110 98 ;
        RECT 97.394 93.133 98 110 ;
        RECT 93.254 97.273 110 98 ;
        RECT 97.348 93.179 98 110 ;
        RECT 93.3 97.227 110 98 ;
        RECT 97.302 93.225 98 110 ;
        RECT 93.346 97.181 110 98 ;
        RECT 97.256 93.271 98 110 ;
        RECT 93.392 97.135 110 98 ;
        RECT 97.21 93.317 98 110 ;
        RECT 93.438 97.089 110 98 ;
        RECT 97.164 93.363 98 110 ;
        RECT 93.484 97.043 110 98 ;
        RECT 97.118 93.409 98 110 ;
        RECT 93.53 96.997 110 98 ;
        RECT 97.072 93.455 98 110 ;
        RECT 93.576 96.951 110 98 ;
        RECT 97.026 93.501 98 110 ;
        RECT 93.622 96.905 110 98 ;
        RECT 96.98 93.547 98 110 ;
        RECT 93.668 96.859 110 98 ;
        RECT 96.934 93.593 98 110 ;
        RECT 93.714 96.813 110 98 ;
        RECT 96.888 93.639 98 110 ;
        RECT 93.76 96.767 110 98 ;
        RECT 96.842 93.685 98 110 ;
        RECT 93.806 96.721 110 98 ;
        RECT 96.796 93.731 98 110 ;
        RECT 93.852 96.675 110 98 ;
        RECT 96.75 93.777 98 110 ;
        RECT 93.898 96.629 110 98 ;
        RECT 96.704 93.823 98 110 ;
        RECT 93.944 96.583 110 98 ;
        RECT 96.658 93.869 98 110 ;
        RECT 93.99 96.537 110 98 ;
        RECT 96.612 93.915 98 110 ;
        RECT 94.036 96.491 110 98 ;
        RECT 96.566 93.961 98 110 ;
        RECT 94.082 96.445 110 98 ;
        RECT 96.52 94.007 98 110 ;
        RECT 94.128 96.399 110 98 ;
        RECT 96.474 94.053 98 110 ;
        RECT 94.174 96.353 110 98 ;
        RECT 96.428 94.099 98 110 ;
        RECT 94.22 96.307 110 98 ;
        RECT 96.382 94.145 98 110 ;
        RECT 94.266 96.261 110 98 ;
        RECT 96.336 94.191 98 110 ;
        RECT 94.312 96.215 110 98 ;
        RECT 96.29 94.237 98 110 ;
        RECT 94.358 96.169 110 98 ;
        RECT 96.244 94.283 98 110 ;
        RECT 94.404 96.123 110 98 ;
        RECT 96.198 94.329 98 110 ;
        RECT 94.45 96.077 110 98 ;
        RECT 96.152 94.375 98 110 ;
        RECT 94.496 96.031 110 98 ;
        RECT 96.106 94.421 98 110 ;
        RECT 94.542 95.985 110 98 ;
        RECT 96.06 94.467 98 110 ;
        RECT 94.588 95.939 110 98 ;
        RECT 96.014 94.513 98 110 ;
        RECT 94.634 95.893 110 98 ;
        RECT 95.968 94.559 98 110 ;
        RECT 94.68 95.847 110 98 ;
        RECT 95.922 94.605 98 110 ;
        RECT 94.726 95.801 110 98 ;
        RECT 95.876 94.651 98 110 ;
        RECT 94.772 95.755 110 98 ;
        RECT 95.83 94.697 98 110 ;
        RECT 94.818 95.709 110 98 ;
        RECT 95.784 94.743 98 110 ;
        RECT 94.864 95.663 110 98 ;
        RECT 95.738 94.789 98 110 ;
        RECT 94.91 95.617 110 98 ;
        RECT 95.692 94.835 98 110 ;
        RECT 94.956 95.571 110 98 ;
        RECT 95.646 94.881 98 110 ;
        RECT 95.002 95.525 110 98 ;
        RECT 95.6 94.927 98 110 ;
        RECT 95.048 95.479 110 98 ;
        RECT 95.554 94.973 98 110 ;
        RECT 95.094 95.433 110 98 ;
        RECT 95.508 95.019 98 110 ;
        RECT 95.14 95.387 110 98 ;
        RECT 95.462 95.065 98 110 ;
        RECT 95.186 95.341 110 98 ;
        RECT 95.416 95.111 98 110 ;
        RECT 95.232 95.295 110 98 ;
        RECT 95.37 95.157 98 110 ;
        RECT 95.278 95.249 110 98 ;
        RECT 95.324 95.203 98 110 ;
      LAYER MET4 ;
        RECT 99.55 91 110 98 ;
        RECT 91 99.527 100.884 99.589 ;
        RECT 91 99.527 100.838 99.635 ;
        RECT 91 99.527 100.792 99.681 ;
        RECT 91 99.527 100.746 99.727 ;
        RECT 91 99.527 100.7 99.773 ;
        RECT 91 99.527 100.654 99.819 ;
        RECT 91 99.527 100.608 99.865 ;
        RECT 91 99.527 100.562 99.911 ;
        RECT 91 99.527 100.516 99.957 ;
        RECT 91 99.527 100.47 100.003 ;
        RECT 91 99.527 100.424 100.049 ;
        RECT 91 99.527 100.378 100.095 ;
        RECT 91 99.527 100.332 100.141 ;
        RECT 91 99.527 100.286 100.187 ;
        RECT 91 99.527 100.24 100.233 ;
        RECT 91 99.527 100.194 100.279 ;
        RECT 91 99.527 100.148 100.325 ;
        RECT 91 99.527 100.102 100.371 ;
        RECT 91 99.527 100.056 100.417 ;
        RECT 91 99.527 100.01 100.463 ;
        RECT 91 99.527 99.964 100.509 ;
        RECT 91 99.527 99.918 100.555 ;
        RECT 91 99.527 99.872 100.601 ;
        RECT 91 99.527 99.826 100.647 ;
        RECT 91 99.527 99.78 100.693 ;
        RECT 91 99.527 99.734 100.739 ;
        RECT 91 99.527 99.688 100.785 ;
        RECT 91 99.527 99.642 100.831 ;
        RECT 91 99.527 99.596 100.877 ;
        RECT 91.046 99.481 100.93 99.543 ;
        RECT 99.518 91.016 99.55 100.916 ;
        RECT 91.092 99.435 100.976 99.497 ;
        RECT 99.472 91.055 99.518 100.955 ;
        RECT 91.138 99.389 101.022 99.451 ;
        RECT 99.426 91.101 99.472 101.001 ;
        RECT 91.184 99.343 101.068 99.405 ;
        RECT 99.38 91.147 99.426 101.047 ;
        RECT 91.23 99.297 101.114 99.359 ;
        RECT 99.334 91.193 99.38 101.093 ;
        RECT 91.276 99.251 101.16 99.313 ;
        RECT 99.288 91.239 99.334 101.139 ;
        RECT 91.322 99.205 101.206 99.267 ;
        RECT 99.242 91.285 99.288 101.185 ;
        RECT 91.368 99.159 101.252 99.221 ;
        RECT 99.196 91.331 99.242 101.231 ;
        RECT 91.414 99.113 101.298 99.175 ;
        RECT 99.15 91.377 99.196 101.277 ;
        RECT 91.46 99.067 101.344 99.129 ;
        RECT 99.104 91.423 99.15 101.323 ;
        RECT 91.506 99.021 101.39 99.083 ;
        RECT 99.058 91.469 99.104 101.369 ;
        RECT 91.552 98.975 101.436 99.037 ;
        RECT 99.012 91.515 99.058 101.415 ;
        RECT 91.598 98.929 101.482 98.991 ;
        RECT 98.966 91.561 99.012 101.461 ;
        RECT 91.644 98.883 101.528 98.945 ;
        RECT 98.92 91.607 98.966 101.507 ;
        RECT 91.69 98.837 101.574 98.899 ;
        RECT 98.874 91.653 98.92 101.553 ;
        RECT 91.736 98.791 101.62 98.853 ;
        RECT 98.828 91.699 98.874 101.599 ;
        RECT 91.782 98.745 101.666 98.807 ;
        RECT 98.782 91.745 98.828 101.645 ;
        RECT 91.828 98.699 101.712 98.761 ;
        RECT 98.736 91.791 98.782 101.691 ;
        RECT 91.874 98.653 101.758 98.715 ;
        RECT 98.69 91.837 98.736 101.737 ;
        RECT 91.92 98.607 101.804 98.669 ;
        RECT 98.644 91.883 98.69 101.783 ;
        RECT 91.966 98.561 101.85 98.623 ;
        RECT 98.598 91.929 98.644 101.829 ;
        RECT 92.012 98.515 101.896 98.577 ;
        RECT 98.552 91.975 98.598 101.875 ;
        RECT 92.058 98.469 101.942 98.531 ;
        RECT 98.506 92.021 98.552 101.921 ;
        RECT 92.104 98.423 101.988 98.485 ;
        RECT 98.46 92.067 98.506 101.967 ;
        RECT 92.15 98.377 102.034 98.439 ;
        RECT 98.414 92.113 98.46 102.013 ;
        RECT 92.196 98.331 102.08 98.393 ;
        RECT 98.368 92.159 98.414 102.059 ;
        RECT 92.242 98.285 102.126 98.347 ;
        RECT 98.322 92.205 98.368 102.105 ;
        RECT 92.288 98.239 102.172 98.301 ;
        RECT 98.276 92.251 98.322 102.151 ;
        RECT 92.334 98.193 102.218 98.255 ;
        RECT 98.23 92.297 98.276 102.197 ;
        RECT 92.38 98.147 102.264 98.209 ;
        RECT 98.184 92.343 98.23 102.243 ;
        RECT 92.426 98.101 102.31 98.163 ;
        RECT 98.138 92.389 98.184 102.289 ;
        RECT 92.472 98.055 102.356 98.117 ;
        RECT 98.092 92.435 98.138 102.335 ;
        RECT 92.518 98.009 102.402 98.071 ;
        RECT 98.046 92.481 98.092 102.381 ;
        RECT 92.564 97.963 102.448 98.024 ;
        RECT 98 92.527 98.046 102.427 ;
        RECT 91 99.527 98 110 ;
        RECT 92.61 97.917 110 98 ;
        RECT 97.992 92.554 98 110 ;
        RECT 92.656 97.871 110 98 ;
        RECT 97.946 92.581 98 110 ;
        RECT 92.702 97.825 110 98 ;
        RECT 97.9 92.627 98 110 ;
        RECT 92.748 97.779 110 98 ;
        RECT 97.854 92.673 98 110 ;
        RECT 92.794 97.733 110 98 ;
        RECT 97.808 92.719 98 110 ;
        RECT 92.84 97.687 110 98 ;
        RECT 97.762 92.765 98 110 ;
        RECT 92.886 97.641 110 98 ;
        RECT 97.716 92.811 98 110 ;
        RECT 92.932 97.595 110 98 ;
        RECT 97.67 92.857 98 110 ;
        RECT 92.978 97.549 110 98 ;
        RECT 97.624 92.903 98 110 ;
        RECT 93.024 97.503 110 98 ;
        RECT 97.578 92.949 98 110 ;
        RECT 93.07 97.457 110 98 ;
        RECT 97.532 92.995 98 110 ;
        RECT 93.116 97.411 110 98 ;
        RECT 97.486 93.041 98 110 ;
        RECT 93.162 97.365 110 98 ;
        RECT 97.44 93.087 98 110 ;
        RECT 93.208 97.319 110 98 ;
        RECT 97.394 93.133 98 110 ;
        RECT 93.254 97.273 110 98 ;
        RECT 97.348 93.179 98 110 ;
        RECT 93.3 97.227 110 98 ;
        RECT 97.302 93.225 98 110 ;
        RECT 93.346 97.181 110 98 ;
        RECT 97.256 93.271 98 110 ;
        RECT 93.392 97.135 110 98 ;
        RECT 97.21 93.317 98 110 ;
        RECT 93.438 97.089 110 98 ;
        RECT 97.164 93.363 98 110 ;
        RECT 93.484 97.043 110 98 ;
        RECT 97.118 93.409 98 110 ;
        RECT 93.53 96.997 110 98 ;
        RECT 97.072 93.455 98 110 ;
        RECT 93.576 96.951 110 98 ;
        RECT 97.026 93.501 98 110 ;
        RECT 93.622 96.905 110 98 ;
        RECT 96.98 93.547 98 110 ;
        RECT 93.668 96.859 110 98 ;
        RECT 96.934 93.593 98 110 ;
        RECT 93.714 96.813 110 98 ;
        RECT 96.888 93.639 98 110 ;
        RECT 93.76 96.767 110 98 ;
        RECT 96.842 93.685 98 110 ;
        RECT 93.806 96.721 110 98 ;
        RECT 96.796 93.731 98 110 ;
        RECT 93.852 96.675 110 98 ;
        RECT 96.75 93.777 98 110 ;
        RECT 93.898 96.629 110 98 ;
        RECT 96.704 93.823 98 110 ;
        RECT 93.944 96.583 110 98 ;
        RECT 96.658 93.869 98 110 ;
        RECT 93.99 96.537 110 98 ;
        RECT 96.612 93.915 98 110 ;
        RECT 94.036 96.491 110 98 ;
        RECT 96.566 93.961 98 110 ;
        RECT 94.082 96.445 110 98 ;
        RECT 96.52 94.007 98 110 ;
        RECT 94.128 96.399 110 98 ;
        RECT 96.474 94.053 98 110 ;
        RECT 94.174 96.353 110 98 ;
        RECT 96.428 94.099 98 110 ;
        RECT 94.22 96.307 110 98 ;
        RECT 96.382 94.145 98 110 ;
        RECT 94.266 96.261 110 98 ;
        RECT 96.336 94.191 98 110 ;
        RECT 94.312 96.215 110 98 ;
        RECT 96.29 94.237 98 110 ;
        RECT 94.358 96.169 110 98 ;
        RECT 96.244 94.283 98 110 ;
        RECT 94.404 96.123 110 98 ;
        RECT 96.198 94.329 98 110 ;
        RECT 94.45 96.077 110 98 ;
        RECT 96.152 94.375 98 110 ;
        RECT 94.496 96.031 110 98 ;
        RECT 96.106 94.421 98 110 ;
        RECT 94.542 95.985 110 98 ;
        RECT 96.06 94.467 98 110 ;
        RECT 94.588 95.939 110 98 ;
        RECT 96.014 94.513 98 110 ;
        RECT 94.634 95.893 110 98 ;
        RECT 95.968 94.559 98 110 ;
        RECT 94.68 95.847 110 98 ;
        RECT 95.922 94.605 98 110 ;
        RECT 94.726 95.801 110 98 ;
        RECT 95.876 94.651 98 110 ;
        RECT 94.772 95.755 110 98 ;
        RECT 95.83 94.697 98 110 ;
        RECT 94.818 95.709 110 98 ;
        RECT 95.784 94.743 98 110 ;
        RECT 94.864 95.663 110 98 ;
        RECT 95.738 94.789 98 110 ;
        RECT 94.91 95.617 110 98 ;
        RECT 95.692 94.835 98 110 ;
        RECT 94.956 95.571 110 98 ;
        RECT 95.646 94.881 98 110 ;
        RECT 95.002 95.525 110 98 ;
        RECT 95.6 94.927 98 110 ;
        RECT 95.048 95.479 110 98 ;
        RECT 95.554 94.973 98 110 ;
        RECT 95.094 95.433 110 98 ;
        RECT 95.508 95.019 98 110 ;
        RECT 95.14 95.387 110 98 ;
        RECT 95.462 95.065 98 110 ;
        RECT 95.186 95.341 110 98 ;
        RECT 95.416 95.111 98 110 ;
        RECT 95.232 95.295 110 98 ;
        RECT 95.37 95.157 98 110 ;
        RECT 95.278 95.249 110 98 ;
        RECT 95.324 95.203 98 110 ;
      LAYER MET3 ;
        RECT 99.55 91 110 98 ;
        RECT 91 99.527 100.884 99.589 ;
        RECT 91 99.527 100.838 99.635 ;
        RECT 91 99.527 100.792 99.681 ;
        RECT 91 99.527 100.746 99.727 ;
        RECT 91 99.527 100.7 99.773 ;
        RECT 91 99.527 100.654 99.819 ;
        RECT 91 99.527 100.608 99.865 ;
        RECT 91 99.527 100.562 99.911 ;
        RECT 91 99.527 100.516 99.957 ;
        RECT 91 99.527 100.47 100.003 ;
        RECT 91 99.527 100.424 100.049 ;
        RECT 91 99.527 100.378 100.095 ;
        RECT 91 99.527 100.332 100.141 ;
        RECT 91 99.527 100.286 100.187 ;
        RECT 91 99.527 100.24 100.233 ;
        RECT 91 99.527 100.194 100.279 ;
        RECT 91 99.527 100.148 100.325 ;
        RECT 91 99.527 100.102 100.371 ;
        RECT 91 99.527 100.056 100.417 ;
        RECT 91 99.527 100.01 100.463 ;
        RECT 91 99.527 99.964 100.509 ;
        RECT 91 99.527 99.918 100.555 ;
        RECT 91 99.527 99.872 100.601 ;
        RECT 91 99.527 99.826 100.647 ;
        RECT 91 99.527 99.78 100.693 ;
        RECT 91 99.527 99.734 100.739 ;
        RECT 91 99.527 99.688 100.785 ;
        RECT 91 99.527 99.642 100.831 ;
        RECT 91 99.527 99.596 100.877 ;
        RECT 91.046 99.481 100.93 99.543 ;
        RECT 99.518 91.016 99.55 100.916 ;
        RECT 91.092 99.435 100.976 99.497 ;
        RECT 99.472 91.055 99.518 100.955 ;
        RECT 91.138 99.389 101.022 99.451 ;
        RECT 99.426 91.101 99.472 101.001 ;
        RECT 91.184 99.343 101.068 99.405 ;
        RECT 99.38 91.147 99.426 101.047 ;
        RECT 91.23 99.297 101.114 99.359 ;
        RECT 99.334 91.193 99.38 101.093 ;
        RECT 91.276 99.251 101.16 99.313 ;
        RECT 99.288 91.239 99.334 101.139 ;
        RECT 91.322 99.205 101.206 99.267 ;
        RECT 99.242 91.285 99.288 101.185 ;
        RECT 91.368 99.159 101.252 99.221 ;
        RECT 99.196 91.331 99.242 101.231 ;
        RECT 91.414 99.113 101.298 99.175 ;
        RECT 99.15 91.377 99.196 101.277 ;
        RECT 91.46 99.067 101.344 99.129 ;
        RECT 99.104 91.423 99.15 101.323 ;
        RECT 91.506 99.021 101.39 99.083 ;
        RECT 99.058 91.469 99.104 101.369 ;
        RECT 91.552 98.975 101.436 99.037 ;
        RECT 99.012 91.515 99.058 101.415 ;
        RECT 91.598 98.929 101.482 98.991 ;
        RECT 98.966 91.561 99.012 101.461 ;
        RECT 91.644 98.883 101.528 98.945 ;
        RECT 98.92 91.607 98.966 101.507 ;
        RECT 91.69 98.837 101.574 98.899 ;
        RECT 98.874 91.653 98.92 101.553 ;
        RECT 91.736 98.791 101.62 98.853 ;
        RECT 98.828 91.699 98.874 101.599 ;
        RECT 91.782 98.745 101.666 98.807 ;
        RECT 98.782 91.745 98.828 101.645 ;
        RECT 91.828 98.699 101.712 98.761 ;
        RECT 98.736 91.791 98.782 101.691 ;
        RECT 91.874 98.653 101.758 98.715 ;
        RECT 98.69 91.837 98.736 101.737 ;
        RECT 91.92 98.607 101.804 98.669 ;
        RECT 98.644 91.883 98.69 101.783 ;
        RECT 91.966 98.561 101.85 98.623 ;
        RECT 98.598 91.929 98.644 101.829 ;
        RECT 92.012 98.515 101.896 98.577 ;
        RECT 98.552 91.975 98.598 101.875 ;
        RECT 92.058 98.469 101.942 98.531 ;
        RECT 98.506 92.021 98.552 101.921 ;
        RECT 92.104 98.423 101.988 98.485 ;
        RECT 98.46 92.067 98.506 101.967 ;
        RECT 92.15 98.377 102.034 98.439 ;
        RECT 98.414 92.113 98.46 102.013 ;
        RECT 92.196 98.331 102.08 98.393 ;
        RECT 98.368 92.159 98.414 102.059 ;
        RECT 92.242 98.285 102.126 98.347 ;
        RECT 98.322 92.205 98.368 102.105 ;
        RECT 92.288 98.239 102.172 98.301 ;
        RECT 98.276 92.251 98.322 102.151 ;
        RECT 92.334 98.193 102.218 98.255 ;
        RECT 98.23 92.297 98.276 102.197 ;
        RECT 92.38 98.147 102.264 98.209 ;
        RECT 98.184 92.343 98.23 102.243 ;
        RECT 92.426 98.101 102.31 98.163 ;
        RECT 98.138 92.389 98.184 102.289 ;
        RECT 92.472 98.055 102.356 98.117 ;
        RECT 98.092 92.435 98.138 102.335 ;
        RECT 92.518 98.009 102.402 98.071 ;
        RECT 98.046 92.481 98.092 102.381 ;
        RECT 92.564 97.963 102.448 98.024 ;
        RECT 98 92.527 98.046 102.427 ;
        RECT 91 99.527 98 110 ;
        RECT 92.61 97.917 110 98 ;
        RECT 97.992 92.554 98 110 ;
        RECT 92.656 97.871 110 98 ;
        RECT 97.946 92.581 98 110 ;
        RECT 92.702 97.825 110 98 ;
        RECT 97.9 92.627 98 110 ;
        RECT 92.748 97.779 110 98 ;
        RECT 97.854 92.673 98 110 ;
        RECT 92.794 97.733 110 98 ;
        RECT 97.808 92.719 98 110 ;
        RECT 92.84 97.687 110 98 ;
        RECT 97.762 92.765 98 110 ;
        RECT 92.886 97.641 110 98 ;
        RECT 97.716 92.811 98 110 ;
        RECT 92.932 97.595 110 98 ;
        RECT 97.67 92.857 98 110 ;
        RECT 92.978 97.549 110 98 ;
        RECT 97.624 92.903 98 110 ;
        RECT 93.024 97.503 110 98 ;
        RECT 97.578 92.949 98 110 ;
        RECT 93.07 97.457 110 98 ;
        RECT 97.532 92.995 98 110 ;
        RECT 93.116 97.411 110 98 ;
        RECT 97.486 93.041 98 110 ;
        RECT 93.162 97.365 110 98 ;
        RECT 97.44 93.087 98 110 ;
        RECT 93.208 97.319 110 98 ;
        RECT 97.394 93.133 98 110 ;
        RECT 93.254 97.273 110 98 ;
        RECT 97.348 93.179 98 110 ;
        RECT 93.3 97.227 110 98 ;
        RECT 97.302 93.225 98 110 ;
        RECT 93.346 97.181 110 98 ;
        RECT 97.256 93.271 98 110 ;
        RECT 93.392 97.135 110 98 ;
        RECT 97.21 93.317 98 110 ;
        RECT 93.438 97.089 110 98 ;
        RECT 97.164 93.363 98 110 ;
        RECT 93.484 97.043 110 98 ;
        RECT 97.118 93.409 98 110 ;
        RECT 93.53 96.997 110 98 ;
        RECT 97.072 93.455 98 110 ;
        RECT 93.576 96.951 110 98 ;
        RECT 97.026 93.501 98 110 ;
        RECT 93.622 96.905 110 98 ;
        RECT 96.98 93.547 98 110 ;
        RECT 93.668 96.859 110 98 ;
        RECT 96.934 93.593 98 110 ;
        RECT 93.714 96.813 110 98 ;
        RECT 96.888 93.639 98 110 ;
        RECT 93.76 96.767 110 98 ;
        RECT 96.842 93.685 98 110 ;
        RECT 93.806 96.721 110 98 ;
        RECT 96.796 93.731 98 110 ;
        RECT 93.852 96.675 110 98 ;
        RECT 96.75 93.777 98 110 ;
        RECT 93.898 96.629 110 98 ;
        RECT 96.704 93.823 98 110 ;
        RECT 93.944 96.583 110 98 ;
        RECT 96.658 93.869 98 110 ;
        RECT 93.99 96.537 110 98 ;
        RECT 96.612 93.915 98 110 ;
        RECT 94.036 96.491 110 98 ;
        RECT 96.566 93.961 98 110 ;
        RECT 94.082 96.445 110 98 ;
        RECT 96.52 94.007 98 110 ;
        RECT 94.128 96.399 110 98 ;
        RECT 96.474 94.053 98 110 ;
        RECT 94.174 96.353 110 98 ;
        RECT 96.428 94.099 98 110 ;
        RECT 94.22 96.307 110 98 ;
        RECT 96.382 94.145 98 110 ;
        RECT 94.266 96.261 110 98 ;
        RECT 96.336 94.191 98 110 ;
        RECT 94.312 96.215 110 98 ;
        RECT 96.29 94.237 98 110 ;
        RECT 94.358 96.169 110 98 ;
        RECT 96.244 94.283 98 110 ;
        RECT 94.404 96.123 110 98 ;
        RECT 96.198 94.329 98 110 ;
        RECT 94.45 96.077 110 98 ;
        RECT 96.152 94.375 98 110 ;
        RECT 94.496 96.031 110 98 ;
        RECT 96.106 94.421 98 110 ;
        RECT 94.542 95.985 110 98 ;
        RECT 96.06 94.467 98 110 ;
        RECT 94.588 95.939 110 98 ;
        RECT 96.014 94.513 98 110 ;
        RECT 94.634 95.893 110 98 ;
        RECT 95.968 94.559 98 110 ;
        RECT 94.68 95.847 110 98 ;
        RECT 95.922 94.605 98 110 ;
        RECT 94.726 95.801 110 98 ;
        RECT 95.876 94.651 98 110 ;
        RECT 94.772 95.755 110 98 ;
        RECT 95.83 94.697 98 110 ;
        RECT 94.818 95.709 110 98 ;
        RECT 95.784 94.743 98 110 ;
        RECT 94.864 95.663 110 98 ;
        RECT 95.738 94.789 98 110 ;
        RECT 94.91 95.617 110 98 ;
        RECT 95.692 94.835 98 110 ;
        RECT 94.956 95.571 110 98 ;
        RECT 95.646 94.881 98 110 ;
        RECT 95.002 95.525 110 98 ;
        RECT 95.6 94.927 98 110 ;
        RECT 95.048 95.479 110 98 ;
        RECT 95.554 94.973 98 110 ;
        RECT 95.094 95.433 110 98 ;
        RECT 95.508 95.019 98 110 ;
        RECT 95.14 95.387 110 98 ;
        RECT 95.462 95.065 98 110 ;
        RECT 95.186 95.341 110 98 ;
        RECT 95.416 95.111 98 110 ;
        RECT 95.232 95.295 110 98 ;
        RECT 95.37 95.157 98 110 ;
        RECT 95.278 95.249 110 98 ;
        RECT 95.324 95.203 98 110 ;
      LAYER MET2 ;
        RECT 99.55 91 110 98 ;
        RECT 91 99.527 100.884 99.589 ;
        RECT 91 99.527 100.838 99.635 ;
        RECT 91 99.527 100.792 99.681 ;
        RECT 91 99.527 100.746 99.727 ;
        RECT 91 99.527 100.7 99.773 ;
        RECT 91 99.527 100.654 99.819 ;
        RECT 91 99.527 100.608 99.865 ;
        RECT 91 99.527 100.562 99.911 ;
        RECT 91 99.527 100.516 99.957 ;
        RECT 91 99.527 100.47 100.003 ;
        RECT 91 99.527 100.424 100.049 ;
        RECT 91 99.527 100.378 100.095 ;
        RECT 91 99.527 100.332 100.141 ;
        RECT 91 99.527 100.286 100.187 ;
        RECT 91 99.527 100.24 100.233 ;
        RECT 91 99.527 100.194 100.279 ;
        RECT 91 99.527 100.148 100.325 ;
        RECT 91 99.527 100.102 100.371 ;
        RECT 91 99.527 100.056 100.417 ;
        RECT 91 99.527 100.01 100.463 ;
        RECT 91 99.527 99.964 100.509 ;
        RECT 91 99.527 99.918 100.555 ;
        RECT 91 99.527 99.872 100.601 ;
        RECT 91 99.527 99.826 100.647 ;
        RECT 91 99.527 99.78 100.693 ;
        RECT 91 99.527 99.734 100.739 ;
        RECT 91 99.527 99.688 100.785 ;
        RECT 91 99.527 99.642 100.831 ;
        RECT 91 99.527 99.596 100.877 ;
        RECT 91.046 99.481 100.93 99.543 ;
        RECT 99.518 91.016 99.55 100.916 ;
        RECT 91.092 99.435 100.976 99.497 ;
        RECT 99.472 91.055 99.518 100.955 ;
        RECT 91.138 99.389 101.022 99.451 ;
        RECT 99.426 91.101 99.472 101.001 ;
        RECT 91.184 99.343 101.068 99.405 ;
        RECT 99.38 91.147 99.426 101.047 ;
        RECT 91.23 99.297 101.114 99.359 ;
        RECT 99.334 91.193 99.38 101.093 ;
        RECT 91.276 99.251 101.16 99.313 ;
        RECT 99.288 91.239 99.334 101.139 ;
        RECT 91.322 99.205 101.206 99.267 ;
        RECT 99.242 91.285 99.288 101.185 ;
        RECT 91.368 99.159 101.252 99.221 ;
        RECT 99.196 91.331 99.242 101.231 ;
        RECT 91.414 99.113 101.298 99.175 ;
        RECT 99.15 91.377 99.196 101.277 ;
        RECT 91.46 99.067 101.344 99.129 ;
        RECT 99.104 91.423 99.15 101.323 ;
        RECT 91.506 99.021 101.39 99.083 ;
        RECT 99.058 91.469 99.104 101.369 ;
        RECT 91.552 98.975 101.436 99.037 ;
        RECT 99.012 91.515 99.058 101.415 ;
        RECT 91.598 98.929 101.482 98.991 ;
        RECT 98.966 91.561 99.012 101.461 ;
        RECT 91.644 98.883 101.528 98.945 ;
        RECT 98.92 91.607 98.966 101.507 ;
        RECT 91.69 98.837 101.574 98.899 ;
        RECT 98.874 91.653 98.92 101.553 ;
        RECT 91.736 98.791 101.62 98.853 ;
        RECT 98.828 91.699 98.874 101.599 ;
        RECT 91.782 98.745 101.666 98.807 ;
        RECT 98.782 91.745 98.828 101.645 ;
        RECT 91.828 98.699 101.712 98.761 ;
        RECT 98.736 91.791 98.782 101.691 ;
        RECT 91.874 98.653 101.758 98.715 ;
        RECT 98.69 91.837 98.736 101.737 ;
        RECT 91.92 98.607 101.804 98.669 ;
        RECT 98.644 91.883 98.69 101.783 ;
        RECT 91.966 98.561 101.85 98.623 ;
        RECT 98.598 91.929 98.644 101.829 ;
        RECT 92.012 98.515 101.896 98.577 ;
        RECT 98.552 91.975 98.598 101.875 ;
        RECT 92.058 98.469 101.942 98.531 ;
        RECT 98.506 92.021 98.552 101.921 ;
        RECT 92.104 98.423 101.988 98.485 ;
        RECT 98.46 92.067 98.506 101.967 ;
        RECT 92.15 98.377 102.034 98.439 ;
        RECT 98.414 92.113 98.46 102.013 ;
        RECT 92.196 98.331 102.08 98.393 ;
        RECT 98.368 92.159 98.414 102.059 ;
        RECT 92.242 98.285 102.126 98.347 ;
        RECT 98.322 92.205 98.368 102.105 ;
        RECT 92.288 98.239 102.172 98.301 ;
        RECT 98.276 92.251 98.322 102.151 ;
        RECT 92.334 98.193 102.218 98.255 ;
        RECT 98.23 92.297 98.276 102.197 ;
        RECT 92.38 98.147 102.264 98.209 ;
        RECT 98.184 92.343 98.23 102.243 ;
        RECT 92.426 98.101 102.31 98.163 ;
        RECT 98.138 92.389 98.184 102.289 ;
        RECT 92.472 98.055 102.356 98.117 ;
        RECT 98.092 92.435 98.138 102.335 ;
        RECT 92.518 98.009 102.402 98.071 ;
        RECT 98.046 92.481 98.092 102.381 ;
        RECT 92.564 97.963 102.448 98.024 ;
        RECT 98 92.527 98.046 102.427 ;
        RECT 91 99.527 98 110 ;
        RECT 92.61 97.917 110 98 ;
        RECT 97.992 92.554 98 110 ;
        RECT 92.656 97.871 110 98 ;
        RECT 97.946 92.581 98 110 ;
        RECT 92.702 97.825 110 98 ;
        RECT 97.9 92.627 98 110 ;
        RECT 92.748 97.779 110 98 ;
        RECT 97.854 92.673 98 110 ;
        RECT 92.794 97.733 110 98 ;
        RECT 97.808 92.719 98 110 ;
        RECT 92.84 97.687 110 98 ;
        RECT 97.762 92.765 98 110 ;
        RECT 92.886 97.641 110 98 ;
        RECT 97.716 92.811 98 110 ;
        RECT 92.932 97.595 110 98 ;
        RECT 97.67 92.857 98 110 ;
        RECT 92.978 97.549 110 98 ;
        RECT 97.624 92.903 98 110 ;
        RECT 93.024 97.503 110 98 ;
        RECT 97.578 92.949 98 110 ;
        RECT 93.07 97.457 110 98 ;
        RECT 97.532 92.995 98 110 ;
        RECT 93.116 97.411 110 98 ;
        RECT 97.486 93.041 98 110 ;
        RECT 93.162 97.365 110 98 ;
        RECT 97.44 93.087 98 110 ;
        RECT 93.208 97.319 110 98 ;
        RECT 97.394 93.133 98 110 ;
        RECT 93.254 97.273 110 98 ;
        RECT 97.348 93.179 98 110 ;
        RECT 93.3 97.227 110 98 ;
        RECT 97.302 93.225 98 110 ;
        RECT 93.346 97.181 110 98 ;
        RECT 97.256 93.271 98 110 ;
        RECT 93.392 97.135 110 98 ;
        RECT 97.21 93.317 98 110 ;
        RECT 93.438 97.089 110 98 ;
        RECT 97.164 93.363 98 110 ;
        RECT 93.484 97.043 110 98 ;
        RECT 97.118 93.409 98 110 ;
        RECT 93.53 96.997 110 98 ;
        RECT 97.072 93.455 98 110 ;
        RECT 93.576 96.951 110 98 ;
        RECT 97.026 93.501 98 110 ;
        RECT 93.622 96.905 110 98 ;
        RECT 96.98 93.547 98 110 ;
        RECT 93.668 96.859 110 98 ;
        RECT 96.934 93.593 98 110 ;
        RECT 93.714 96.813 110 98 ;
        RECT 96.888 93.639 98 110 ;
        RECT 93.76 96.767 110 98 ;
        RECT 96.842 93.685 98 110 ;
        RECT 93.806 96.721 110 98 ;
        RECT 96.796 93.731 98 110 ;
        RECT 93.852 96.675 110 98 ;
        RECT 96.75 93.777 98 110 ;
        RECT 93.898 96.629 110 98 ;
        RECT 96.704 93.823 98 110 ;
        RECT 93.944 96.583 110 98 ;
        RECT 96.658 93.869 98 110 ;
        RECT 93.99 96.537 110 98 ;
        RECT 96.612 93.915 98 110 ;
        RECT 94.036 96.491 110 98 ;
        RECT 96.566 93.961 98 110 ;
        RECT 94.082 96.445 110 98 ;
        RECT 96.52 94.007 98 110 ;
        RECT 94.128 96.399 110 98 ;
        RECT 96.474 94.053 98 110 ;
        RECT 94.174 96.353 110 98 ;
        RECT 96.428 94.099 98 110 ;
        RECT 94.22 96.307 110 98 ;
        RECT 96.382 94.145 98 110 ;
        RECT 94.266 96.261 110 98 ;
        RECT 96.336 94.191 98 110 ;
        RECT 94.312 96.215 110 98 ;
        RECT 96.29 94.237 98 110 ;
        RECT 94.358 96.169 110 98 ;
        RECT 96.244 94.283 98 110 ;
        RECT 94.404 96.123 110 98 ;
        RECT 96.198 94.329 98 110 ;
        RECT 94.45 96.077 110 98 ;
        RECT 96.152 94.375 98 110 ;
        RECT 94.496 96.031 110 98 ;
        RECT 96.106 94.421 98 110 ;
        RECT 94.542 95.985 110 98 ;
        RECT 96.06 94.467 98 110 ;
        RECT 94.588 95.939 110 98 ;
        RECT 96.014 94.513 98 110 ;
        RECT 94.634 95.893 110 98 ;
        RECT 95.968 94.559 98 110 ;
        RECT 94.68 95.847 110 98 ;
        RECT 95.922 94.605 98 110 ;
        RECT 94.726 95.801 110 98 ;
        RECT 95.876 94.651 98 110 ;
        RECT 94.772 95.755 110 98 ;
        RECT 95.83 94.697 98 110 ;
        RECT 94.818 95.709 110 98 ;
        RECT 95.784 94.743 98 110 ;
        RECT 94.864 95.663 110 98 ;
        RECT 95.738 94.789 98 110 ;
        RECT 94.91 95.617 110 98 ;
        RECT 95.692 94.835 98 110 ;
        RECT 94.956 95.571 110 98 ;
        RECT 95.646 94.881 98 110 ;
        RECT 95.002 95.525 110 98 ;
        RECT 95.6 94.927 98 110 ;
        RECT 95.048 95.479 110 98 ;
        RECT 95.554 94.973 98 110 ;
        RECT 95.094 95.433 110 98 ;
        RECT 95.508 95.019 98 110 ;
        RECT 95.14 95.387 110 98 ;
        RECT 95.462 95.065 98 110 ;
        RECT 95.186 95.341 110 98 ;
        RECT 95.416 95.111 98 110 ;
        RECT 95.232 95.295 110 98 ;
        RECT 95.37 95.157 98 110 ;
        RECT 95.278 95.249 110 98 ;
        RECT 95.324 95.203 98 110 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.016941 LAYER MET4 ;
    ANTENNAPARTIALMETALAREA 0.016941 LAYER MET3 ;
    ANTENNAPARTIALMETALAREA 0.016941 LAYER MET2 ;
    ANTENNAPARTIALCUTAREA 17.6256 LAYER VIA4 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 29.16 LAYER VIA2 ;
    PORT
      LAYER MET5 ;
        RECT 28.316 51.426 45.238 51.515 ;
        RECT 28.27 51.472 45.192 51.561 ;
        RECT 28.224 51.518 45.146 51.607 ;
        RECT 28.178 51.564 45.1 51.653 ;
        RECT 28.132 51.61 45.054 51.699 ;
        RECT 28.086 51.656 45.008 51.745 ;
        RECT 28.04 51.702 44.962 51.791 ;
        RECT 27.994 51.748 44.916 51.837 ;
        RECT 27.948 51.794 44.87 51.883 ;
        RECT 27.902 51.84 44.824 51.929 ;
        RECT 27.856 51.886 44.778 51.975 ;
        RECT 27.81 51.932 44.732 52.021 ;
        RECT 27.764 51.978 44.686 52.067 ;
        RECT 27.718 52.024 44.64 52.113 ;
        RECT 27.672 52.07 44.594 52.159 ;
        RECT 27.626 52.116 44.548 52.205 ;
        RECT 27.58 52.162 44.502 52.251 ;
        RECT 27.534 52.208 44.456 52.297 ;
        RECT 27.488 52.254 44.41 52.343 ;
        RECT 27.442 52.3 44.364 52.389 ;
        RECT 27.396 52.346 44.318 52.435 ;
        RECT 27.35 52.392 44.272 52.481 ;
        RECT 27.304 52.438 44.226 52.527 ;
        RECT 27.258 52.484 44.18 52.573 ;
        RECT 27.212 52.53 44.134 52.619 ;
        RECT 27.166 52.576 44.088 52.665 ;
        RECT 27.12 52.622 44.042 52.711 ;
        RECT 27.074 52.668 43.996 52.757 ;
        RECT 27.028 52.714 43.95 52.803 ;
        RECT 26.982 52.76 43.904 52.849 ;
        RECT 26.936 52.806 43.858 52.895 ;
        RECT 26.89 52.852 43.812 52.941 ;
        RECT 26.844 52.898 43.766 52.987 ;
        RECT 26.798 52.944 43.72 53.033 ;
        RECT 26.752 52.99 43.674 53.079 ;
        RECT 26.706 53.036 43.628 53.125 ;
        RECT 26.66 53.082 43.582 53.171 ;
        RECT 26.614 53.128 43.536 53.217 ;
        RECT 26.568 53.174 43.49 53.263 ;
        RECT 26.522 53.22 43.444 53.309 ;
        RECT 26.476 53.266 43.398 53.355 ;
        RECT 26.43 53.312 43.352 53.401 ;
        RECT 26.384 53.358 43.306 53.447 ;
        RECT 26.338 53.404 43.26 53.493 ;
        RECT 26.292 53.45 43.214 53.539 ;
        RECT 26.246 53.496 43.168 53.585 ;
        RECT 26.2 53.542 43.122 53.631 ;
        RECT 26.154 53.588 43.076 53.677 ;
        RECT 26.108 53.634 43.03 53.723 ;
        RECT 26.062 53.68 42.984 53.769 ;
        RECT 26.016 53.726 42.938 53.815 ;
        RECT 25.97 53.772 42.892 53.861 ;
        RECT 25.924 53.818 42.846 53.907 ;
        RECT 25.878 53.864 42.8 53.953 ;
        RECT 25.832 53.91 42.754 53.999 ;
        RECT 25.786 53.956 42.708 54.045 ;
        RECT 25.74 54.002 42.662 54.091 ;
        RECT 25.694 54.048 42.616 54.137 ;
        RECT 25.648 54.094 42.57 54.183 ;
        RECT 25.602 54.14 42.524 54.229 ;
        RECT 25.556 54.186 42.478 54.275 ;
        RECT 25.51 54.232 42.432 54.321 ;
        RECT 25.464 54.278 42.386 54.367 ;
        RECT 25.418 54.324 42.34 54.413 ;
        RECT 25.372 54.37 42.294 54.459 ;
        RECT 25.326 54.416 42.248 54.505 ;
        RECT 25.28 54.462 42.202 54.551 ;
        RECT 25.234 54.508 42.156 54.597 ;
        RECT 25.188 54.554 42.11 54.643 ;
        RECT 25.142 54.6 42.064 54.689 ;
        RECT 25.096 54.646 42.018 54.735 ;
        RECT 25.05 54.692 41.972 54.781 ;
        RECT 25.004 54.738 41.926 54.827 ;
        RECT 24.958 54.784 41.88 54.873 ;
        RECT 24.912 54.83 41.834 54.919 ;
        RECT 24.866 54.876 41.788 54.965 ;
        RECT 24.82 54.922 41.742 55.011 ;
        RECT 24.774 54.968 41.696 55.057 ;
        RECT 24.728 55.014 41.65 55.103 ;
        RECT 24.682 55.06 41.604 55.149 ;
        RECT 24.636 55.106 41.558 55.195 ;
        RECT 24.59 55.152 41.512 55.241 ;
        RECT 24.544 55.198 41.466 55.287 ;
        RECT 24.498 55.244 41.42 55.333 ;
        RECT 24.452 55.29 41.374 55.379 ;
        RECT 24.406 55.336 41.328 55.425 ;
        RECT 24.36 55.382 41.282 55.471 ;
        RECT 24.314 55.428 41.236 55.517 ;
        RECT 24.268 55.474 41.19 55.563 ;
        RECT 24.222 55.52 41.144 55.609 ;
        RECT 24.176 55.566 41.098 55.655 ;
        RECT 24.13 55.612 41.052 55.701 ;
        RECT 24.084 55.658 41.006 55.747 ;
        RECT 24.038 55.704 40.96 55.793 ;
        RECT 23.992 55.75 40.914 55.839 ;
        RECT 23.946 55.796 40.868 55.885 ;
        RECT 23.9 55.842 40.822 55.931 ;
        RECT 23.854 55.888 40.776 55.977 ;
        RECT 23.808 55.934 40.73 56.023 ;
        RECT 23.762 55.98 40.684 56.069 ;
        RECT 23.716 56.026 40.638 56.115 ;
        RECT 23.67 56.072 40.592 56.161 ;
        RECT 23.624 56.118 40.546 56.207 ;
        RECT 23.578 56.164 40.5 56.253 ;
        RECT 23.532 56.21 40.454 56.299 ;
        RECT 23.486 56.256 40.408 56.345 ;
        RECT 23.44 56.302 40.362 56.391 ;
        RECT 23.394 56.348 40.316 56.437 ;
        RECT 23.348 56.394 40.27 56.483 ;
        RECT 23.302 56.44 40.224 56.529 ;
        RECT 23.256 56.486 40.178 56.575 ;
        RECT 23.21 56.532 40.132 56.621 ;
        RECT 23.164 56.578 40.086 56.667 ;
        RECT 23.118 56.624 40.04 56.713 ;
        RECT 23.072 56.67 39.994 56.759 ;
        RECT 23.026 56.716 39.948 56.805 ;
        RECT 22.98 56.762 39.902 56.851 ;
        RECT 22.934 56.808 39.856 56.897 ;
        RECT 22.888 56.854 39.81 56.943 ;
        RECT 22.842 56.9 39.764 56.989 ;
        RECT 22.796 56.946 39.718 57.035 ;
        RECT 22.75 56.992 39.672 57.081 ;
        RECT 22.704 57.038 39.626 57.127 ;
        RECT 22.658 57.084 39.58 57.173 ;
        RECT 22.612 57.13 39.534 57.219 ;
        RECT 22.566 57.176 39.488 57.265 ;
        RECT 22.52 57.222 39.442 57.311 ;
        RECT 22.474 57.268 39.396 57.357 ;
        RECT 22.428 57.314 39.35 57.403 ;
        RECT 22.382 57.36 39.304 57.449 ;
        RECT 22.336 57.406 39.258 57.495 ;
        RECT 22.29 57.452 39.212 57.541 ;
        RECT 22.244 57.498 39.166 57.587 ;
        RECT 22.198 57.544 39.12 57.633 ;
        RECT 22.152 57.59 39.074 57.679 ;
        RECT 22.106 57.636 39.028 57.725 ;
        RECT 22.06 57.682 38.982 57.771 ;
        RECT 22.014 57.728 38.936 57.817 ;
        RECT 21.968 57.774 38.89 57.863 ;
        RECT 21.922 57.82 38.844 57.909 ;
        RECT 21.876 57.866 38.798 57.955 ;
        RECT 21.83 57.912 38.752 58.001 ;
        RECT 21.784 57.958 38.706 58.047 ;
        RECT 21.738 58.004 38.66 58.093 ;
        RECT 21.692 58.05 38.614 58.139 ;
        RECT 21.646 58.096 38.568 58.185 ;
        RECT 21.6 58.142 38.522 58.231 ;
        RECT 21.554 58.188 38.476 58.277 ;
        RECT 21.508 58.234 38.43 58.323 ;
        RECT 21.462 58.28 38.384 58.369 ;
        RECT 21.416 58.326 38.338 58.415 ;
        RECT 21.37 58.372 38.292 58.461 ;
        RECT 21.324 58.418 38.246 58.507 ;
        RECT 21.278 58.464 38.2 58.553 ;
        RECT 21.232 58.51 38.154 58.599 ;
        RECT 21.186 58.556 38.108 58.645 ;
        RECT 21.14 58.602 38.062 58.691 ;
        RECT 21.094 58.648 38.016 58.737 ;
        RECT 21.048 58.694 37.97 58.783 ;
        RECT 21.002 58.74 37.924 58.829 ;
        RECT 20.956 58.786 37.878 58.875 ;
        RECT 20.91 58.832 37.832 58.921 ;
        RECT 20.864 58.878 37.786 58.967 ;
        RECT 20.818 58.924 37.74 59.013 ;
        RECT 20.772 58.97 37.694 59.059 ;
        RECT 20.726 59.016 37.648 59.105 ;
        RECT 20.68 59.062 37.602 59.151 ;
        RECT 20.634 59.108 37.556 59.197 ;
        RECT 20.588 59.154 37.51 59.243 ;
        RECT 20.542 59.2 37.464 59.289 ;
        RECT 20.496 59.246 37.418 59.335 ;
        RECT 20.45 59.292 37.372 59.381 ;
        RECT 20.404 59.338 37.326 59.427 ;
        RECT 20.358 59.384 37.28 59.473 ;
        RECT 20.312 59.43 37.234 59.519 ;
        RECT 20.266 59.476 37.188 59.565 ;
        RECT 20.22 59.522 37.142 59.611 ;
        RECT 20.174 59.568 37.096 59.657 ;
        RECT 20.128 59.614 37.05 59.703 ;
        RECT 20.082 59.66 37.004 59.749 ;
        RECT 20.036 59.706 36.958 59.795 ;
        RECT 19.99 59.752 36.912 59.841 ;
        RECT 19.944 59.798 36.866 59.887 ;
        RECT 19.898 59.844 36.82 59.933 ;
        RECT 19.852 59.89 36.774 59.979 ;
        RECT 19.806 59.936 36.728 60.025 ;
        RECT 19.76 59.982 36.682 60.071 ;
        RECT 19.714 60.028 36.636 60.117 ;
        RECT 19.668 60.074 36.59 60.163 ;
        RECT 19.622 60.12 36.544 60.209 ;
        RECT 19.576 60.166 36.498 60.255 ;
        RECT 19.53 60.212 36.452 60.301 ;
        RECT 19.484 60.258 36.406 60.347 ;
        RECT 19.438 60.304 36.36 60.393 ;
        RECT 19.392 60.35 36.314 60.439 ;
        RECT 19.346 60.396 36.268 60.485 ;
        RECT 19.3 60.442 36.222 60.531 ;
        RECT 19.254 60.488 36.176 60.577 ;
        RECT 19.208 60.534 36.13 60.623 ;
        RECT 19.162 60.58 36.084 60.669 ;
        RECT 19.116 60.626 36.038 60.715 ;
        RECT 19.07 60.672 35.992 60.761 ;
        RECT 19.024 60.718 35.946 60.807 ;
        RECT 18.978 60.764 35.9 60.853 ;
        RECT 18.932 60.81 35.854 60.899 ;
        RECT 18.886 60.856 35.808 60.945 ;
        RECT 18.84 60.902 35.762 60.991 ;
        RECT 18.794 60.948 35.716 61.037 ;
        RECT 18.748 60.994 35.67 61.083 ;
        RECT 18.702 61.04 35.624 61.129 ;
        RECT 18.656 61.086 35.578 61.175 ;
        RECT 18.61 61.132 35.532 61.221 ;
        RECT 18.564 61.178 35.486 61.267 ;
        RECT 18.518 61.224 35.44 61.313 ;
        RECT 18.472 61.27 35.394 61.359 ;
        RECT 18.426 61.316 35.348 61.405 ;
        RECT 18.38 61.362 35.302 61.451 ;
        RECT 18.334 61.408 35.256 61.497 ;
        RECT 18.288 61.454 35.21 61.543 ;
        RECT 18.242 61.5 35.164 61.589 ;
        RECT 18.196 61.546 35.118 61.635 ;
        RECT 18.15 61.592 35.072 61.681 ;
        RECT 18.104 61.638 35.026 61.727 ;
        RECT 18.058 61.684 34.98 61.773 ;
        RECT 18.012 61.73 34.934 61.819 ;
        RECT 17.966 61.776 34.888 61.865 ;
        RECT 17.92 61.822 34.842 61.911 ;
        RECT 17.874 61.868 34.796 61.957 ;
        RECT 17.828 61.914 34.75 62.003 ;
        RECT 17.782 61.96 34.704 62.049 ;
        RECT 17.736 62.006 34.658 62.095 ;
        RECT 17.69 62.052 34.612 62.141 ;
        RECT 17.644 62.098 34.566 62.187 ;
        RECT 17.598 62.144 34.52 62.233 ;
        RECT 17.552 62.19 34.474 62.279 ;
        RECT 17.506 62.236 34.428 62.325 ;
        RECT 17.46 62.282 34.382 62.371 ;
        RECT 17.414 62.328 34.336 62.417 ;
        RECT 17.368 62.374 34.29 62.463 ;
        RECT 17.322 62.42 34.244 62.509 ;
        RECT 17.276 62.466 34.198 62.555 ;
        RECT 17.23 62.512 34.152 62.601 ;
        RECT 17.184 62.558 34.106 62.647 ;
        RECT 17.138 62.604 34.06 62.693 ;
        RECT 17.092 62.65 34.014 62.739 ;
        RECT 17.046 62.696 33.968 62.785 ;
        RECT 17 62.742 33.922 62.831 ;
        RECT 17 62.742 33.876 62.877 ;
        RECT 17 62.742 33.83 62.923 ;
        RECT 17 62.742 33.784 62.969 ;
        RECT 17 62.742 33.738 63.015 ;
        RECT 17 62.742 33.692 63.061 ;
        RECT 17 62.742 33.646 63.107 ;
        RECT 17 62.742 33.6 63.153 ;
        RECT 17 62.742 33.554 63.199 ;
        RECT 17 62.742 33.508 63.245 ;
        RECT 17 62.742 33.462 63.291 ;
        RECT 17 62.742 33.416 63.337 ;
        RECT 17 62.742 33.37 63.383 ;
        RECT 17 62.742 33.324 63.429 ;
        RECT 17 62.742 33.278 63.475 ;
        RECT 17 62.742 33.232 63.521 ;
        RECT 17 62.742 33.186 63.567 ;
        RECT 17 62.742 33.14 63.613 ;
        RECT 17 62.742 33.094 63.659 ;
        RECT 17 62.742 33.048 63.705 ;
        RECT 17 62.742 33.002 63.751 ;
        RECT 17 62.742 32.956 63.797 ;
        RECT 17 62.742 32.91 63.843 ;
        RECT 17 62.742 32.864 63.889 ;
        RECT 17 62.742 32.818 63.935 ;
        RECT 17 62.742 32.772 63.981 ;
        RECT 17 62.742 32.726 64.027 ;
        RECT 17 62.742 32.68 64.073 ;
        RECT 17 62.742 32.634 64.119 ;
        RECT 17 62.742 32.588 64.165 ;
        RECT 17 62.742 32.542 64.211 ;
        RECT 17 62.742 32.496 64.257 ;
        RECT 17 62.742 32.45 64.303 ;
        RECT 17 62.742 32.404 64.349 ;
        RECT 17 62.742 32.358 64.395 ;
        RECT 17 62.742 32.312 64.441 ;
        RECT 17 62.742 32.266 64.487 ;
        RECT 17 62.742 32.22 64.533 ;
        RECT 17 62.742 32.174 64.579 ;
        RECT 17 62.742 32.128 64.625 ;
        RECT 17 62.742 32.082 64.671 ;
        RECT 17 62.742 32.036 64.717 ;
        RECT 17 62.742 31.99 64.763 ;
        RECT 17 62.742 31.944 64.809 ;
        RECT 17 62.742 31.898 64.855 ;
        RECT 17 62.742 31.852 64.901 ;
        RECT 17 62.742 31.806 64.947 ;
        RECT 17 62.742 31.76 64.993 ;
        RECT 17 62.742 31.714 65.039 ;
        RECT 17 62.742 31.668 65.085 ;
        RECT 17 62.742 31.622 65.131 ;
        RECT 17 62.742 31.576 65.177 ;
        RECT 17 62.742 31.53 65.223 ;
        RECT 17 62.742 31.484 65.269 ;
        RECT 17 62.742 31.438 65.315 ;
        RECT 17 62.742 31.392 65.361 ;
        RECT 17 62.742 31.346 65.407 ;
        RECT 17 62.742 31.3 65.453 ;
        RECT 17 62.742 31.254 65.499 ;
        RECT 17 62.742 31.208 65.545 ;
        RECT 17 62.742 31.162 65.591 ;
        RECT 17 62.742 31.116 65.637 ;
        RECT 17 62.742 31.07 65.683 ;
        RECT 17 62.742 31.024 65.729 ;
        RECT 17 62.742 30.978 65.775 ;
        RECT 17 62.742 30.932 65.821 ;
        RECT 17 62.742 30.886 65.867 ;
        RECT 17 62.742 30.84 65.913 ;
        RECT 17 62.742 30.794 65.959 ;
        RECT 17 62.742 30.748 66.005 ;
        RECT 17 62.742 30.702 66.051 ;
        RECT 17 62.742 30.656 66.097 ;
        RECT 17 62.742 30.61 66.143 ;
        RECT 17 62.742 30.564 66.189 ;
        RECT 17 62.742 30.518 66.235 ;
        RECT 17 62.742 30.472 66.281 ;
        RECT 17 62.742 30.426 66.327 ;
        RECT 17 62.742 30.38 66.373 ;
        RECT 17 62.742 30.334 66.419 ;
        RECT 17 62.742 30.288 66.465 ;
        RECT 17 62.742 30.242 66.511 ;
        RECT 17 62.742 30.196 66.557 ;
        RECT 17 62.742 30.15 66.603 ;
        RECT 17 62.742 30.104 66.649 ;
        RECT 17 62.742 30.058 66.695 ;
        RECT 17 62.742 30.012 66.741 ;
        RECT 17 62.742 29.966 66.787 ;
        RECT 17 62.742 29.92 66.833 ;
        RECT 17 62.742 29.874 66.879 ;
        RECT 17 62.742 29.828 66.925 ;
        RECT 17 62.742 29.782 66.971 ;
        RECT 17 62.742 29.736 67.017 ;
        RECT 17 62.742 29.69 67.063 ;
        RECT 17 62.742 29.644 67.109 ;
        RECT 17 62.742 29.598 67.155 ;
        RECT 17 62.742 29.552 67.201 ;
        RECT 17 62.742 29.506 67.247 ;
        RECT 17 62.742 29.46 67.293 ;
        RECT 17 62.742 29.414 67.339 ;
        RECT 17 62.742 29.368 67.385 ;
        RECT 17 62.742 29.322 67.431 ;
        RECT 17 62.742 29.276 67.477 ;
        RECT 17 62.742 29.23 67.523 ;
        RECT 17 62.742 29.184 67.569 ;
        RECT 17 62.742 29.138 67.615 ;
        RECT 17 62.742 29.092 67.661 ;
        RECT 17 62.742 29.046 67.707 ;
        RECT 17 62.742 29 110 ;
        RECT 92.47 78.5 110 89.5 ;
        RECT 78.5 92.447 94.034 92.509 ;
        RECT 78.5 92.447 93.988 92.555 ;
        RECT 78.5 92.447 93.942 92.601 ;
        RECT 78.5 92.447 93.896 92.647 ;
        RECT 78.5 92.447 93.85 92.693 ;
        RECT 78.5 92.447 93.804 92.739 ;
        RECT 78.5 92.447 93.758 92.785 ;
        RECT 78.5 92.447 93.712 92.831 ;
        RECT 78.5 92.447 93.666 92.877 ;
        RECT 78.5 92.447 93.62 92.923 ;
        RECT 78.5 92.447 93.574 92.969 ;
        RECT 78.5 92.447 93.528 93.015 ;
        RECT 78.5 92.447 93.482 93.061 ;
        RECT 78.5 92.447 93.436 93.107 ;
        RECT 78.5 92.447 93.39 93.153 ;
        RECT 78.5 92.447 93.344 93.199 ;
        RECT 78.5 92.447 93.298 93.245 ;
        RECT 78.5 92.447 93.252 93.291 ;
        RECT 78.5 92.447 93.206 93.337 ;
        RECT 78.5 92.447 93.16 93.383 ;
        RECT 78.5 92.447 93.114 93.429 ;
        RECT 78.5 92.447 93.068 93.475 ;
        RECT 78.5 92.447 93.022 93.521 ;
        RECT 78.5 92.447 92.976 93.567 ;
        RECT 78.5 92.447 92.93 93.613 ;
        RECT 78.5 92.447 92.884 93.659 ;
        RECT 78.5 92.447 92.838 93.705 ;
        RECT 78.5 92.447 92.792 93.751 ;
        RECT 78.5 92.447 92.746 93.797 ;
        RECT 78.5 92.447 92.7 93.843 ;
        RECT 78.5 92.447 92.654 93.889 ;
        RECT 78.5 92.447 92.608 93.935 ;
        RECT 78.5 92.447 92.562 93.981 ;
        RECT 78.5 92.447 92.516 94.027 ;
        RECT 78.546 92.401 94.08 92.463 ;
        RECT 92.444 78.513 92.47 94.063 ;
        RECT 78.592 92.355 94.126 92.417 ;
        RECT 92.398 78.549 92.444 94.099 ;
        RECT 78.638 92.309 94.172 92.371 ;
        RECT 92.352 78.595 92.398 94.145 ;
        RECT 78.684 92.263 94.218 92.325 ;
        RECT 92.306 78.641 92.352 94.191 ;
        RECT 78.73 92.217 94.264 92.279 ;
        RECT 92.26 78.687 92.306 94.237 ;
        RECT 78.776 92.171 94.31 92.233 ;
        RECT 92.214 78.733 92.26 94.283 ;
        RECT 78.822 92.125 94.356 92.187 ;
        RECT 92.168 78.779 92.214 94.329 ;
        RECT 78.868 92.079 94.402 92.141 ;
        RECT 92.122 78.825 92.168 94.375 ;
        RECT 78.914 92.033 94.448 92.095 ;
        RECT 92.076 78.871 92.122 94.421 ;
        RECT 78.96 91.987 94.494 92.049 ;
        RECT 92.03 78.917 92.076 94.467 ;
        RECT 79.006 91.941 94.54 92.003 ;
        RECT 91.984 78.963 92.03 94.513 ;
        RECT 79.052 91.895 94.586 91.957 ;
        RECT 91.938 79.009 91.984 94.559 ;
        RECT 79.098 91.849 94.632 91.911 ;
        RECT 91.892 79.055 91.938 94.605 ;
        RECT 79.144 91.803 94.678 91.865 ;
        RECT 91.846 79.101 91.892 94.651 ;
        RECT 79.19 91.757 94.724 91.819 ;
        RECT 91.8 79.147 91.846 94.697 ;
        RECT 79.236 91.711 94.77 91.773 ;
        RECT 91.754 79.193 91.8 94.743 ;
        RECT 79.282 91.665 94.816 91.727 ;
        RECT 91.708 79.239 91.754 94.789 ;
        RECT 79.328 91.619 94.862 91.681 ;
        RECT 91.662 79.285 91.708 94.835 ;
        RECT 79.374 91.573 94.908 91.635 ;
        RECT 91.616 79.331 91.662 94.881 ;
        RECT 79.42 91.527 94.954 91.589 ;
        RECT 91.57 79.377 91.616 94.927 ;
        RECT 79.466 91.481 95 91.543 ;
        RECT 91.524 79.423 91.57 94.973 ;
        RECT 79.512 91.435 95.046 91.497 ;
        RECT 91.478 79.469 91.524 95.019 ;
        RECT 79.558 91.389 95.092 91.451 ;
        RECT 91.432 79.515 91.478 95.065 ;
        RECT 79.604 91.343 95.138 91.405 ;
        RECT 91.386 79.561 91.432 95.111 ;
        RECT 79.65 91.297 95.184 91.359 ;
        RECT 91.34 79.607 91.386 95.157 ;
        RECT 79.696 91.251 95.23 91.313 ;
        RECT 91.294 79.653 91.34 95.203 ;
        RECT 79.742 91.205 95.276 91.267 ;
        RECT 91.248 79.699 91.294 95.249 ;
        RECT 79.788 91.159 95.322 91.221 ;
        RECT 91.202 79.745 91.248 95.295 ;
        RECT 79.834 91.113 95.368 91.175 ;
        RECT 91.156 79.791 91.202 95.341 ;
        RECT 79.88 91.067 95.414 91.129 ;
        RECT 91.11 79.837 91.156 95.387 ;
        RECT 79.926 91.021 95.46 91.083 ;
        RECT 91.064 79.883 91.11 95.433 ;
        RECT 79.972 90.975 95.506 91.037 ;
        RECT 91.018 79.929 91.064 95.479 ;
        RECT 80.018 90.929 95.552 90.991 ;
        RECT 90.972 79.975 91.018 95.525 ;
        RECT 80.064 90.883 95.598 90.945 ;
        RECT 90.926 80.021 90.972 95.571 ;
        RECT 80.11 90.837 95.644 90.899 ;
        RECT 90.88 80.067 90.926 95.617 ;
        RECT 80.156 90.791 95.69 90.853 ;
        RECT 90.834 80.113 90.88 95.663 ;
        RECT 80.202 90.745 95.736 90.807 ;
        RECT 90.788 80.159 90.834 95.709 ;
        RECT 80.248 90.699 95.782 90.761 ;
        RECT 90.742 80.205 90.788 95.755 ;
        RECT 80.294 90.653 95.828 90.715 ;
        RECT 90.696 80.251 90.742 95.801 ;
        RECT 80.34 90.607 95.874 90.669 ;
        RECT 90.65 80.297 90.696 95.847 ;
        RECT 80.386 90.561 95.92 90.623 ;
        RECT 90.604 80.343 90.65 95.893 ;
        RECT 80.432 90.515 95.966 90.577 ;
        RECT 90.558 80.389 90.604 95.939 ;
        RECT 80.478 90.469 96.012 90.531 ;
        RECT 90.512 80.435 90.558 95.985 ;
        RECT 80.524 90.423 96.058 90.485 ;
        RECT 90.466 80.481 90.512 96.031 ;
        RECT 80.57 90.377 96.104 90.439 ;
        RECT 90.42 80.527 90.466 96.077 ;
        RECT 80.616 90.331 96.15 90.393 ;
        RECT 90.374 80.573 90.42 96.123 ;
        RECT 80.662 90.285 96.196 90.347 ;
        RECT 90.328 80.619 90.374 96.169 ;
        RECT 80.708 90.239 96.242 90.301 ;
        RECT 90.282 80.665 90.328 96.215 ;
        RECT 80.754 90.193 96.288 90.255 ;
        RECT 90.236 80.711 90.282 96.261 ;
        RECT 80.8 90.147 96.334 90.209 ;
        RECT 90.19 80.757 90.236 96.307 ;
        RECT 80.846 90.101 96.38 90.163 ;
        RECT 90.144 80.803 90.19 96.353 ;
        RECT 80.892 90.055 96.426 90.117 ;
        RECT 90.098 80.849 90.144 96.399 ;
        RECT 80.938 90.009 96.472 90.071 ;
        RECT 90.052 80.895 90.098 96.445 ;
        RECT 80.984 89.963 96.518 90.025 ;
        RECT 90.006 80.941 90.052 96.491 ;
        RECT 81.03 89.917 96.564 89.979 ;
        RECT 89.96 80.987 90.006 96.537 ;
        RECT 81.076 89.871 96.61 89.933 ;
        RECT 89.914 81.033 89.96 96.583 ;
        RECT 81.122 89.825 96.656 89.887 ;
        RECT 89.868 81.079 89.914 96.629 ;
        RECT 81.168 89.779 96.702 89.841 ;
        RECT 89.822 81.125 89.868 96.675 ;
        RECT 81.214 89.733 96.748 89.795 ;
        RECT 89.776 81.171 89.822 96.721 ;
        RECT 81.26 89.687 96.794 89.749 ;
        RECT 89.73 81.217 89.776 96.767 ;
        RECT 81.306 89.641 96.84 89.703 ;
        RECT 89.684 81.263 89.73 96.813 ;
        RECT 81.352 89.595 96.886 89.657 ;
        RECT 89.638 81.309 89.684 96.859 ;
        RECT 81.398 89.549 96.932 89.611 ;
        RECT 89.592 81.355 89.638 96.905 ;
        RECT 81.444 89.503 96.978 89.565 ;
        RECT 89.546 81.401 89.592 96.951 ;
        RECT 81.49 89.457 97.02 89.521 ;
        RECT 89.5 81.447 89.546 96.997 ;
        RECT 78.5 92.447 89.5 110 ;
        RECT 81.536 89.411 110 89.5 ;
        RECT 89.494 81.473 89.5 110 ;
        RECT 81.582 89.365 110 89.5 ;
        RECT 89.448 81.499 89.5 110 ;
        RECT 81.628 89.319 110 89.5 ;
        RECT 89.402 81.545 89.5 110 ;
        RECT 81.674 89.273 110 89.5 ;
        RECT 89.356 81.591 89.5 110 ;
        RECT 81.72 89.227 110 89.5 ;
        RECT 89.31 81.637 89.5 110 ;
        RECT 81.766 89.181 110 89.5 ;
        RECT 89.264 81.683 89.5 110 ;
        RECT 81.812 89.135 110 89.5 ;
        RECT 89.218 81.729 89.5 110 ;
        RECT 81.858 89.089 110 89.5 ;
        RECT 89.172 81.775 89.5 110 ;
        RECT 81.904 89.043 110 89.5 ;
        RECT 89.126 81.821 89.5 110 ;
        RECT 81.95 88.997 110 89.5 ;
        RECT 89.08 81.867 89.5 110 ;
        RECT 81.996 88.951 110 89.5 ;
        RECT 89.034 81.913 89.5 110 ;
        RECT 82.042 88.905 110 89.5 ;
        RECT 88.988 81.959 89.5 110 ;
        RECT 82.088 88.859 110 89.5 ;
        RECT 88.942 82.005 89.5 110 ;
        RECT 82.134 88.813 110 89.5 ;
        RECT 88.896 82.051 89.5 110 ;
        RECT 82.18 88.767 110 89.5 ;
        RECT 88.85 82.097 89.5 110 ;
        RECT 82.226 88.721 110 89.5 ;
        RECT 88.804 82.143 89.5 110 ;
        RECT 82.272 88.675 110 89.5 ;
        RECT 88.758 82.189 89.5 110 ;
        RECT 82.318 88.629 110 89.5 ;
        RECT 88.712 82.235 89.5 110 ;
        RECT 82.364 88.583 110 89.5 ;
        RECT 88.666 82.281 89.5 110 ;
        RECT 82.41 88.537 110 89.5 ;
        RECT 88.62 82.327 89.5 110 ;
        RECT 82.456 88.491 110 89.5 ;
        RECT 88.574 82.373 89.5 110 ;
        RECT 82.502 88.445 110 89.5 ;
        RECT 88.528 82.419 89.5 110 ;
        RECT 82.548 88.399 110 89.5 ;
        RECT 88.482 82.465 89.5 110 ;
        RECT 82.594 88.353 110 89.5 ;
        RECT 88.436 82.511 89.5 110 ;
        RECT 82.64 88.307 110 89.5 ;
        RECT 88.39 82.557 89.5 110 ;
        RECT 82.686 88.261 110 89.5 ;
        RECT 88.344 82.603 89.5 110 ;
        RECT 82.732 88.215 110 89.5 ;
        RECT 88.298 82.649 89.5 110 ;
        RECT 82.778 88.169 110 89.5 ;
        RECT 88.252 82.695 89.5 110 ;
        RECT 82.824 88.123 110 89.5 ;
        RECT 88.206 82.741 89.5 110 ;
        RECT 82.87 88.077 110 89.5 ;
        RECT 88.16 82.787 89.5 110 ;
        RECT 82.916 88.031 110 89.5 ;
        RECT 88.114 82.833 89.5 110 ;
        RECT 82.962 87.985 110 89.5 ;
        RECT 88.068 82.879 89.5 110 ;
        RECT 83.008 87.939 110 89.5 ;
        RECT 88.022 82.925 89.5 110 ;
        RECT 83.054 87.893 110 89.5 ;
        RECT 87.976 82.971 89.5 110 ;
        RECT 83.1 87.847 110 89.5 ;
        RECT 87.93 83.017 89.5 110 ;
        RECT 83.146 87.801 110 89.5 ;
        RECT 87.884 83.063 89.5 110 ;
        RECT 83.192 87.755 110 89.5 ;
        RECT 87.838 83.109 89.5 110 ;
        RECT 83.238 87.709 110 89.5 ;
        RECT 87.792 83.155 89.5 110 ;
        RECT 83.284 87.663 110 89.5 ;
        RECT 87.746 83.201 89.5 110 ;
        RECT 83.33 87.617 110 89.5 ;
        RECT 87.7 83.247 89.5 110 ;
        RECT 83.376 87.571 110 89.5 ;
        RECT 87.654 83.293 89.5 110 ;
        RECT 83.422 87.525 110 89.5 ;
        RECT 87.608 83.339 89.5 110 ;
        RECT 83.468 87.479 110 89.5 ;
        RECT 87.562 83.385 89.5 110 ;
        RECT 83.514 87.433 110 89.5 ;
        RECT 87.516 83.431 89.5 110 ;
        RECT 83.56 87.387 110 89.5 ;
        RECT 87.47 83.477 89.5 110 ;
        RECT 83.606 87.341 110 89.5 ;
        RECT 87.424 83.523 89.5 110 ;
        RECT 83.652 87.295 110 89.5 ;
        RECT 87.378 83.569 89.5 110 ;
        RECT 83.698 87.249 110 89.5 ;
        RECT 87.332 83.615 89.5 110 ;
        RECT 83.744 87.203 110 89.5 ;
        RECT 87.286 83.661 89.5 110 ;
        RECT 83.79 87.157 110 89.5 ;
        RECT 87.24 83.707 89.5 110 ;
        RECT 83.836 87.111 110 89.5 ;
        RECT 87.194 83.753 89.5 110 ;
        RECT 83.882 87.065 110 89.5 ;
        RECT 87.148 83.799 89.5 110 ;
        RECT 83.928 87.019 110 89.5 ;
        RECT 87.102 83.845 89.5 110 ;
        RECT 83.974 86.973 110 89.5 ;
        RECT 87.056 83.891 89.5 110 ;
        RECT 84.02 86.927 110 89.5 ;
        RECT 87.01 83.937 89.5 110 ;
        RECT 84.066 86.881 110 89.5 ;
        RECT 86.964 83.983 89.5 110 ;
        RECT 84.112 86.835 110 89.5 ;
        RECT 86.918 84.029 89.5 110 ;
        RECT 84.158 86.789 110 89.5 ;
        RECT 86.872 84.075 89.5 110 ;
        RECT 84.204 86.743 110 89.5 ;
        RECT 86.826 84.121 89.5 110 ;
        RECT 84.25 86.697 110 89.5 ;
        RECT 86.78 84.167 89.5 110 ;
        RECT 84.296 86.651 110 89.5 ;
        RECT 86.734 84.213 89.5 110 ;
        RECT 84.342 86.605 110 89.5 ;
        RECT 86.688 84.259 89.5 110 ;
        RECT 84.388 86.559 110 89.5 ;
        RECT 86.642 84.305 89.5 110 ;
        RECT 84.434 86.513 110 89.5 ;
        RECT 86.596 84.351 89.5 110 ;
        RECT 84.48 86.467 110 89.5 ;
        RECT 86.55 84.397 89.5 110 ;
        RECT 84.526 86.421 110 89.5 ;
        RECT 86.504 84.443 89.5 110 ;
        RECT 84.572 86.375 110 89.5 ;
        RECT 86.458 84.489 89.5 110 ;
        RECT 84.618 86.329 110 89.5 ;
        RECT 86.412 84.535 89.5 110 ;
        RECT 84.664 86.283 110 89.5 ;
        RECT 86.366 84.581 89.5 110 ;
        RECT 84.71 86.237 110 89.5 ;
        RECT 86.32 84.627 89.5 110 ;
        RECT 84.756 86.191 110 89.5 ;
        RECT 86.274 84.673 89.5 110 ;
        RECT 84.802 86.145 110 89.5 ;
        RECT 86.228 84.719 89.5 110 ;
        RECT 84.848 86.099 110 89.5 ;
        RECT 86.182 84.765 89.5 110 ;
        RECT 84.894 86.053 110 89.5 ;
        RECT 86.136 84.811 89.5 110 ;
        RECT 84.94 86.007 110 89.5 ;
        RECT 86.09 84.857 89.5 110 ;
        RECT 84.986 85.961 110 89.5 ;
        RECT 86.044 84.903 89.5 110 ;
        RECT 85.032 85.915 110 89.5 ;
        RECT 85.998 84.949 89.5 110 ;
        RECT 85.078 85.869 110 89.5 ;
        RECT 85.952 84.995 89.5 110 ;
        RECT 85.124 85.823 110 89.5 ;
        RECT 85.906 85.041 89.5 110 ;
        RECT 85.17 85.777 110 89.5 ;
        RECT 85.86 85.087 89.5 110 ;
        RECT 85.216 85.731 110 89.5 ;
        RECT 85.814 85.133 89.5 110 ;
        RECT 85.262 85.685 110 89.5 ;
        RECT 85.768 85.179 89.5 110 ;
        RECT 85.308 85.639 110 89.5 ;
        RECT 85.722 85.225 89.5 110 ;
        RECT 85.354 85.593 110 89.5 ;
        RECT 85.676 85.271 89.5 110 ;
        RECT 85.4 85.547 110 89.5 ;
        RECT 85.63 85.317 89.5 110 ;
        RECT 85.446 85.501 110 89.5 ;
        RECT 85.584 85.363 89.5 110 ;
        RECT 85.492 85.455 110 89.5 ;
        RECT 85.538 85.409 89.5 110 ;
        RECT 10.032 49.46 26.954 49.549 ;
        RECT 9.986 49.506 26.908 49.595 ;
        RECT 9.94 49.552 26.862 49.641 ;
        RECT 9.894 49.598 26.816 49.687 ;
        RECT 9.848 49.644 26.77 49.733 ;
        RECT 9.802 49.69 26.724 49.779 ;
        RECT 9.756 49.736 26.678 49.825 ;
        RECT 9.71 49.782 26.632 49.871 ;
        RECT 9.664 49.828 26.586 49.917 ;
        RECT 9.618 49.874 26.54 49.963 ;
        RECT 9.572 49.92 26.494 50.009 ;
        RECT 9.526 49.966 26.448 50.055 ;
        RECT 9.48 50.012 26.402 50.101 ;
        RECT 9.434 50.058 26.356 50.147 ;
        RECT 9.388 50.104 26.31 50.193 ;
        RECT 9.342 50.15 26.264 50.239 ;
        RECT 9.296 50.196 26.218 50.285 ;
        RECT 9.25 50.242 26.172 50.331 ;
        RECT 9.204 50.288 26.126 50.377 ;
        RECT 9.158 50.334 26.08 50.423 ;
        RECT 9.112 50.38 26.034 50.469 ;
        RECT 9.066 50.426 25.988 50.515 ;
        RECT 9.02 50.472 25.942 50.561 ;
        RECT 8.974 50.518 25.896 50.607 ;
        RECT 8.928 50.564 25.85 50.653 ;
        RECT 8.882 50.61 25.804 50.699 ;
        RECT 8.836 50.656 25.758 50.745 ;
        RECT 8.79 50.702 25.712 50.791 ;
        RECT 8.744 50.748 25.666 50.837 ;
        RECT 8.698 50.794 25.62 50.883 ;
        RECT 8.652 50.84 25.574 50.929 ;
        RECT 8.606 50.886 25.528 50.975 ;
        RECT 8.56 50.932 25.482 51.021 ;
        RECT 8.514 50.978 25.436 51.067 ;
        RECT 8.468 51.024 25.39 51.113 ;
        RECT 8.422 51.07 25.344 51.159 ;
        RECT 8.376 51.116 25.298 51.205 ;
        RECT 8.33 51.162 25.252 51.251 ;
        RECT 8.284 51.208 25.206 51.297 ;
        RECT 8.238 51.254 25.16 51.343 ;
        RECT 8.192 51.3 25.114 51.389 ;
        RECT 8.146 51.346 25.068 51.435 ;
        RECT 8.1 51.392 25.022 51.481 ;
        RECT 8.054 51.438 24.976 51.527 ;
        RECT 8.008 51.484 24.93 51.573 ;
        RECT 7.962 51.53 24.884 51.619 ;
        RECT 7.916 51.576 24.838 51.665 ;
        RECT 7.87 51.622 24.792 51.711 ;
        RECT 7.824 51.668 24.746 51.757 ;
        RECT 7.778 51.714 24.7 51.803 ;
        RECT 7.732 51.76 24.654 51.849 ;
        RECT 7.686 51.806 24.608 51.895 ;
        RECT 7.64 51.852 24.562 51.941 ;
        RECT 7.594 51.898 24.516 51.987 ;
        RECT 7.548 51.944 24.47 52.033 ;
        RECT 7.502 51.99 24.424 52.079 ;
        RECT 7.456 52.036 24.378 52.125 ;
        RECT 7.41 52.082 24.332 52.171 ;
        RECT 7.364 52.128 24.286 52.217 ;
        RECT 7.318 52.174 24.24 52.263 ;
        RECT 7.272 52.22 24.194 52.309 ;
        RECT 7.226 52.266 24.148 52.355 ;
        RECT 7.18 52.312 24.102 52.401 ;
        RECT 7.134 52.358 24.056 52.447 ;
        RECT 7.088 52.404 24.01 52.493 ;
        RECT 7.042 52.45 23.964 52.539 ;
        RECT 6.996 52.496 23.918 52.585 ;
        RECT 6.95 52.542 23.872 52.631 ;
        RECT 6.904 52.588 23.826 52.677 ;
        RECT 6.858 52.634 23.78 52.723 ;
        RECT 6.812 52.68 23.734 52.769 ;
        RECT 6.766 52.726 23.688 52.815 ;
        RECT 6.72 52.772 23.642 52.861 ;
        RECT 6.674 52.818 23.596 52.907 ;
        RECT 6.628 52.864 23.55 52.953 ;
        RECT 6.582 52.91 23.504 52.999 ;
        RECT 6.536 52.956 23.458 53.045 ;
        RECT 6.49 53.002 23.412 53.091 ;
        RECT 6.444 53.048 23.366 53.137 ;
        RECT 6.398 53.094 23.32 53.183 ;
        RECT 6.352 53.14 23.274 53.229 ;
        RECT 6.306 53.186 23.228 53.275 ;
        RECT 6.26 53.232 23.182 53.321 ;
        RECT 6.214 53.278 23.136 53.367 ;
        RECT 6.168 53.324 23.09 53.413 ;
        RECT 6.122 53.37 23.044 53.459 ;
        RECT 6.076 53.416 22.998 53.505 ;
        RECT 6.03 53.462 22.952 53.551 ;
        RECT 5.984 53.508 22.906 53.597 ;
        RECT 5.938 53.554 22.86 53.643 ;
        RECT 5.892 53.6 22.814 53.689 ;
        RECT 5.846 53.646 22.768 53.735 ;
        RECT 5.8 53.692 22.722 53.781 ;
        RECT 5.754 53.738 22.676 53.827 ;
        RECT 5.708 53.784 22.63 53.873 ;
        RECT 5.662 53.83 22.584 53.919 ;
        RECT 5.616 53.876 22.538 53.965 ;
        RECT 5.57 53.922 22.492 54.011 ;
        RECT 5.524 53.968 22.446 54.057 ;
        RECT 5.478 54.014 22.4 54.103 ;
        RECT 5.432 54.06 22.354 54.149 ;
        RECT 5.386 54.106 22.308 54.195 ;
        RECT 5.34 54.152 22.262 54.241 ;
        RECT 5.294 54.198 22.216 54.287 ;
        RECT 5.248 54.244 22.17 54.333 ;
        RECT 5.202 54.29 22.124 54.379 ;
        RECT 5.156 54.336 22.078 54.425 ;
        RECT 5.11 54.382 22.032 54.471 ;
        RECT 5.064 54.428 21.986 54.517 ;
        RECT 5.018 54.474 21.94 54.563 ;
        RECT 4.972 54.52 21.894 54.609 ;
        RECT 4.926 54.566 21.848 54.655 ;
        RECT 4.88 54.612 21.802 54.701 ;
        RECT 4.834 54.658 21.756 54.747 ;
        RECT 4.788 54.704 21.71 54.793 ;
        RECT 4.742 54.75 21.664 54.839 ;
        RECT 4.696 54.796 21.618 54.885 ;
        RECT 4.65 54.842 21.572 54.931 ;
        RECT 4.604 54.888 21.526 54.977 ;
        RECT 4.558 54.934 21.48 55.023 ;
        RECT 4.512 54.98 21.434 55.069 ;
        RECT 4.466 55.026 21.388 55.115 ;
        RECT 4.42 55.072 21.342 55.161 ;
        RECT 4.374 55.118 21.296 55.207 ;
        RECT 4.328 55.164 21.25 55.253 ;
        RECT 4.282 55.21 21.204 55.299 ;
        RECT 4.236 55.256 21.158 55.345 ;
        RECT 4.19 55.302 21.112 55.391 ;
        RECT 4.144 55.348 21.066 55.437 ;
        RECT 4.098 55.394 21.02 55.483 ;
        RECT 4.052 55.44 20.974 55.529 ;
        RECT 4.006 55.486 20.928 55.575 ;
        RECT 3.96 55.532 20.882 55.621 ;
        RECT 3.914 55.578 20.836 55.667 ;
        RECT 3.868 55.624 20.79 55.713 ;
        RECT 3.822 55.67 20.744 55.759 ;
        RECT 3.776 55.716 20.698 55.805 ;
        RECT 3.73 55.762 20.652 55.851 ;
        RECT 3.684 55.808 20.606 55.897 ;
        RECT 3.638 55.854 20.56 55.943 ;
        RECT 3.592 55.9 20.514 55.989 ;
        RECT 3.546 55.946 20.468 56.035 ;
        RECT 3.5 55.992 20.422 56.081 ;
        RECT 3.5 55.992 20.376 56.127 ;
        RECT 3.5 55.992 20.33 56.173 ;
        RECT 3.5 55.992 20.284 56.219 ;
        RECT 3.5 55.992 20.238 56.265 ;
        RECT 3.5 55.992 20.192 56.311 ;
        RECT 3.5 55.992 20.146 56.357 ;
        RECT 3.5 55.992 20.1 56.403 ;
        RECT 3.5 55.992 20.054 56.449 ;
        RECT 3.5 55.992 20.008 56.495 ;
        RECT 3.5 55.992 19.962 56.541 ;
        RECT 3.5 55.992 19.916 56.587 ;
        RECT 3.5 55.992 19.87 56.633 ;
        RECT 3.5 55.992 19.824 56.679 ;
        RECT 3.5 55.992 19.778 56.725 ;
        RECT 3.5 55.992 19.732 56.771 ;
        RECT 3.5 55.992 19.686 56.817 ;
        RECT 3.5 55.992 19.64 56.863 ;
        RECT 3.5 55.992 19.594 56.909 ;
        RECT 3.5 55.992 19.548 56.955 ;
        RECT 3.5 55.992 19.502 57.001 ;
        RECT 3.5 55.992 19.456 57.047 ;
        RECT 3.5 55.992 19.41 57.093 ;
        RECT 3.5 55.992 19.364 57.139 ;
        RECT 3.5 55.992 19.318 57.185 ;
        RECT 3.5 55.992 19.272 57.231 ;
        RECT 3.5 55.992 19.226 57.277 ;
        RECT 3.5 55.992 19.18 57.323 ;
        RECT 3.5 55.992 19.134 57.369 ;
        RECT 3.5 55.992 19.088 57.415 ;
        RECT 3.5 55.992 19.042 57.461 ;
        RECT 3.5 55.992 18.996 57.507 ;
        RECT 3.5 55.992 18.95 57.553 ;
        RECT 3.5 55.992 18.904 57.599 ;
        RECT 3.5 55.992 18.858 57.645 ;
        RECT 3.5 55.992 18.812 57.691 ;
        RECT 3.5 55.992 18.766 57.737 ;
        RECT 3.5 55.992 18.72 57.783 ;
        RECT 3.5 55.992 18.674 57.829 ;
        RECT 3.5 55.992 18.628 57.875 ;
        RECT 3.5 55.992 18.582 57.921 ;
        RECT 3.5 55.992 18.536 57.967 ;
        RECT 3.5 55.992 18.49 58.013 ;
        RECT 3.5 55.992 18.444 58.059 ;
        RECT 3.5 55.992 18.398 58.105 ;
        RECT 3.5 55.992 18.352 58.151 ;
        RECT 3.5 55.992 18.306 58.197 ;
        RECT 3.5 55.992 18.26 58.243 ;
        RECT 3.5 55.992 18.214 58.289 ;
        RECT 3.5 55.992 18.168 58.335 ;
        RECT 3.5 55.992 18.122 58.381 ;
        RECT 3.5 55.992 18.076 58.427 ;
        RECT 3.5 55.992 18.03 58.473 ;
        RECT 3.5 55.992 17.984 58.519 ;
        RECT 3.5 55.992 17.938 58.565 ;
        RECT 3.5 55.992 17.892 58.611 ;
        RECT 3.5 55.992 17.846 58.657 ;
        RECT 3.5 55.992 17.8 58.703 ;
        RECT 3.5 55.992 17.754 58.749 ;
        RECT 3.5 55.992 17.708 58.795 ;
        RECT 3.5 55.992 17.662 58.841 ;
        RECT 3.5 55.992 17.616 58.887 ;
        RECT 3.5 55.992 17.57 58.933 ;
        RECT 3.5 55.992 17.524 58.979 ;
        RECT 3.5 55.992 17.478 59.025 ;
        RECT 3.5 55.992 17.432 59.071 ;
        RECT 3.5 55.992 17.386 59.117 ;
        RECT 3.5 55.992 17.34 59.163 ;
        RECT 3.5 55.992 17.294 59.209 ;
        RECT 3.5 55.992 17.248 59.255 ;
        RECT 3.5 55.992 17.202 59.301 ;
        RECT 3.5 55.992 17.156 59.347 ;
        RECT 3.5 55.992 17.11 59.393 ;
        RECT 3.5 55.992 17.064 59.439 ;
        RECT 3.5 55.992 17.018 59.485 ;
        RECT 3.5 55.992 16.972 59.531 ;
        RECT 3.5 55.992 16.926 59.577 ;
        RECT 3.5 55.992 16.88 59.623 ;
        RECT 3.5 55.992 16.834 59.669 ;
        RECT 3.5 55.992 16.788 59.715 ;
        RECT 3.5 55.992 16.742 59.761 ;
        RECT 3.5 55.992 16.696 59.807 ;
        RECT 3.5 55.992 16.65 59.853 ;
        RECT 3.5 55.992 16.604 59.899 ;
        RECT 3.5 55.992 16.558 59.945 ;
        RECT 3.5 55.992 16.512 59.991 ;
        RECT 3.5 55.992 16.466 60.037 ;
        RECT 3.5 55.992 16.42 60.083 ;
        RECT 3.5 55.992 16.374 60.129 ;
        RECT 3.5 55.992 16.328 60.175 ;
        RECT 3.5 55.992 16.282 60.221 ;
        RECT 3.5 55.992 16.236 60.267 ;
        RECT 3.5 55.992 16.19 60.313 ;
        RECT 3.5 55.992 16.144 60.359 ;
        RECT 3.5 55.992 16.098 60.405 ;
        RECT 3.5 55.992 16.052 60.451 ;
        RECT 3.5 55.992 16.006 60.497 ;
        RECT 3.5 55.992 15.96 60.543 ;
        RECT 3.5 55.992 15.914 60.589 ;
        RECT 3.5 55.992 15.868 60.635 ;
        RECT 3.5 55.992 15.822 60.681 ;
        RECT 3.5 55.992 15.776 60.727 ;
        RECT 3.5 55.992 15.73 60.773 ;
        RECT 3.5 55.992 15.684 60.819 ;
        RECT 3.5 55.992 15.638 60.865 ;
        RECT 3.5 55.992 15.592 60.911 ;
        RECT 3.5 55.992 15.546 60.957 ;
        RECT 3.5 55.992 15.5 110 ;
        RECT 62.764 17 110 29 ;
        RECT 50.758 28.984 67.73 29.022 ;
        RECT 45.836 33.906 62.765 33.966 ;
        RECT 62.718 17.024 62.764 33.989 ;
        RECT 45.79 33.952 62.718 34.035 ;
        RECT 45.882 33.86 62.811 33.942 ;
        RECT 62.672 17.07 62.718 34.035 ;
        RECT 45.744 33.998 62.672 34.081 ;
        RECT 45.928 33.814 62.857 33.896 ;
        RECT 62.626 17.116 62.672 34.081 ;
        RECT 45.698 34.044 62.626 34.127 ;
        RECT 45.974 33.768 62.903 33.85 ;
        RECT 62.58 17.162 62.626 34.127 ;
        RECT 45.652 34.09 62.58 34.173 ;
        RECT 46.02 33.722 62.949 33.804 ;
        RECT 62.534 17.208 62.58 34.173 ;
        RECT 45.606 34.136 62.534 34.219 ;
        RECT 46.066 33.676 62.995 33.758 ;
        RECT 62.488 17.254 62.534 34.219 ;
        RECT 45.56 34.182 62.488 34.265 ;
        RECT 46.112 33.63 63.041 33.712 ;
        RECT 62.442 17.3 62.488 34.265 ;
        RECT 45.514 34.228 62.442 34.311 ;
        RECT 46.158 33.584 63.087 33.666 ;
        RECT 62.396 17.346 62.442 34.311 ;
        RECT 45.468 34.274 62.396 34.357 ;
        RECT 46.204 33.538 63.133 33.62 ;
        RECT 62.35 17.392 62.396 34.357 ;
        RECT 45.422 34.32 62.35 34.403 ;
        RECT 46.25 33.492 63.179 33.574 ;
        RECT 62.304 17.438 62.35 34.403 ;
        RECT 45.376 34.366 62.304 34.449 ;
        RECT 46.296 33.446 63.225 33.528 ;
        RECT 62.258 17.484 62.304 34.449 ;
        RECT 45.33 34.412 62.258 34.495 ;
        RECT 46.342 33.4 63.271 33.482 ;
        RECT 62.212 17.53 62.258 34.495 ;
        RECT 45.284 34.458 62.212 34.541 ;
        RECT 46.388 33.354 63.317 33.436 ;
        RECT 62.166 17.576 62.212 34.541 ;
        RECT 45.238 34.504 62.166 34.587 ;
        RECT 46.434 33.308 63.363 33.39 ;
        RECT 62.12 17.622 62.166 34.587 ;
        RECT 45.192 34.55 62.12 34.633 ;
        RECT 46.48 33.262 63.409 33.344 ;
        RECT 62.074 17.668 62.12 34.633 ;
        RECT 45.146 34.596 62.074 34.679 ;
        RECT 46.526 33.216 63.455 33.298 ;
        RECT 62.028 17.714 62.074 34.679 ;
        RECT 45.1 34.642 62.028 34.725 ;
        RECT 46.572 33.17 63.501 33.252 ;
        RECT 61.982 17.76 62.028 34.725 ;
        RECT 45.054 34.688 61.982 34.771 ;
        RECT 46.618 33.124 63.547 33.206 ;
        RECT 61.936 17.806 61.982 34.771 ;
        RECT 45.008 34.734 61.936 34.817 ;
        RECT 46.664 33.078 63.593 33.16 ;
        RECT 61.89 17.852 61.936 34.817 ;
        RECT 44.962 34.78 61.89 34.863 ;
        RECT 46.71 33.032 63.639 33.114 ;
        RECT 61.844 17.898 61.89 34.863 ;
        RECT 44.916 34.826 61.844 34.909 ;
        RECT 46.756 32.986 63.685 33.068 ;
        RECT 61.798 17.944 61.844 34.909 ;
        RECT 44.87 34.872 61.798 34.955 ;
        RECT 46.802 32.94 63.731 33.022 ;
        RECT 61.752 17.99 61.798 34.955 ;
        RECT 44.824 34.918 61.752 35.001 ;
        RECT 46.848 32.894 63.777 32.976 ;
        RECT 61.706 18.036 61.752 35.001 ;
        RECT 44.778 34.964 61.706 35.047 ;
        RECT 46.894 32.848 63.823 32.93 ;
        RECT 61.66 18.082 61.706 35.047 ;
        RECT 44.732 35.01 61.66 35.093 ;
        RECT 46.94 32.802 63.869 32.884 ;
        RECT 61.614 18.128 61.66 35.093 ;
        RECT 44.686 35.056 61.614 35.139 ;
        RECT 46.986 32.756 63.915 32.838 ;
        RECT 61.568 18.174 61.614 35.139 ;
        RECT 44.64 35.102 61.568 35.185 ;
        RECT 47.032 32.71 63.961 32.792 ;
        RECT 61.522 18.22 61.568 35.185 ;
        RECT 44.594 35.148 61.522 35.231 ;
        RECT 47.078 32.664 64.007 32.746 ;
        RECT 61.476 18.266 61.522 35.231 ;
        RECT 44.548 35.194 61.476 35.277 ;
        RECT 47.124 32.618 64.053 32.7 ;
        RECT 61.43 18.312 61.476 35.277 ;
        RECT 44.502 35.24 61.43 35.323 ;
        RECT 47.17 32.572 64.099 32.654 ;
        RECT 61.384 18.358 61.43 35.323 ;
        RECT 44.456 35.286 61.384 35.369 ;
        RECT 47.216 32.526 64.145 32.608 ;
        RECT 61.338 18.404 61.384 35.369 ;
        RECT 44.41 35.332 61.338 35.415 ;
        RECT 47.262 32.48 64.191 32.562 ;
        RECT 61.292 18.45 61.338 35.415 ;
        RECT 44.364 35.378 61.292 35.461 ;
        RECT 47.308 32.434 64.237 32.516 ;
        RECT 61.246 18.496 61.292 35.461 ;
        RECT 44.318 35.424 61.246 35.507 ;
        RECT 47.354 32.388 64.283 32.47 ;
        RECT 61.2 18.542 61.246 35.507 ;
        RECT 44.272 35.47 61.2 35.553 ;
        RECT 47.4 32.342 64.329 32.424 ;
        RECT 61.154 18.588 61.2 35.553 ;
        RECT 44.226 35.516 61.154 35.599 ;
        RECT 47.446 32.296 64.375 32.378 ;
        RECT 61.108 18.634 61.154 35.599 ;
        RECT 44.18 35.562 61.108 35.645 ;
        RECT 47.492 32.25 64.421 32.332 ;
        RECT 61.062 18.68 61.108 35.645 ;
        RECT 44.134 35.608 61.062 35.691 ;
        RECT 47.538 32.204 64.467 32.286 ;
        RECT 61.016 18.726 61.062 35.691 ;
        RECT 44.088 35.654 61.016 35.737 ;
        RECT 47.584 32.158 64.513 32.24 ;
        RECT 60.97 18.772 61.016 35.737 ;
        RECT 44.042 35.7 60.97 35.783 ;
        RECT 47.63 32.112 64.559 32.194 ;
        RECT 60.924 18.818 60.97 35.783 ;
        RECT 43.996 35.746 60.924 35.829 ;
        RECT 47.676 32.066 64.605 32.148 ;
        RECT 60.878 18.864 60.924 35.829 ;
        RECT 43.95 35.792 60.878 35.875 ;
        RECT 47.722 32.02 64.651 32.102 ;
        RECT 60.832 18.91 60.878 35.875 ;
        RECT 43.904 35.838 60.832 35.921 ;
        RECT 47.768 31.974 64.697 32.056 ;
        RECT 60.786 18.956 60.832 35.921 ;
        RECT 43.858 35.884 60.786 35.967 ;
        RECT 47.814 31.928 64.743 32.01 ;
        RECT 60.74 19.002 60.786 35.967 ;
        RECT 43.812 35.93 60.74 36.013 ;
        RECT 47.86 31.882 64.789 31.964 ;
        RECT 60.694 19.048 60.74 36.013 ;
        RECT 43.766 35.976 60.694 36.059 ;
        RECT 47.906 31.836 64.835 31.918 ;
        RECT 60.648 19.094 60.694 36.059 ;
        RECT 43.72 36.022 60.648 36.105 ;
        RECT 47.952 31.79 64.881 31.872 ;
        RECT 60.602 19.14 60.648 36.105 ;
        RECT 43.674 36.068 60.602 36.151 ;
        RECT 47.998 31.744 64.927 31.826 ;
        RECT 60.556 19.186 60.602 36.151 ;
        RECT 43.628 36.114 60.556 36.197 ;
        RECT 48.044 31.698 64.973 31.78 ;
        RECT 60.51 19.232 60.556 36.197 ;
        RECT 43.582 36.16 60.51 36.243 ;
        RECT 48.09 31.652 65.019 31.734 ;
        RECT 60.464 19.278 60.51 36.243 ;
        RECT 43.536 36.206 60.464 36.289 ;
        RECT 48.136 31.606 65.065 31.688 ;
        RECT 60.418 19.324 60.464 36.289 ;
        RECT 43.49 36.252 60.418 36.335 ;
        RECT 48.182 31.56 65.111 31.642 ;
        RECT 60.372 19.37 60.418 36.335 ;
        RECT 43.444 36.298 60.372 36.381 ;
        RECT 48.228 31.514 65.157 31.596 ;
        RECT 60.326 19.416 60.372 36.381 ;
        RECT 43.398 36.344 60.326 36.427 ;
        RECT 48.274 31.468 65.203 31.55 ;
        RECT 60.28 19.462 60.326 36.427 ;
        RECT 43.352 36.39 60.28 36.473 ;
        RECT 48.32 31.422 65.249 31.504 ;
        RECT 60.234 19.508 60.28 36.473 ;
        RECT 43.306 36.436 60.234 36.519 ;
        RECT 48.366 31.376 65.295 31.458 ;
        RECT 60.188 19.554 60.234 36.519 ;
        RECT 43.26 36.482 60.188 36.565 ;
        RECT 48.412 31.33 65.341 31.412 ;
        RECT 60.142 19.6 60.188 36.565 ;
        RECT 43.214 36.528 60.142 36.611 ;
        RECT 48.458 31.284 65.387 31.366 ;
        RECT 60.096 19.646 60.142 36.611 ;
        RECT 43.168 36.574 60.096 36.657 ;
        RECT 48.504 31.238 65.433 31.32 ;
        RECT 60.05 19.692 60.096 36.657 ;
        RECT 43.122 36.62 60.05 36.703 ;
        RECT 48.55 31.192 65.479 31.274 ;
        RECT 60.004 19.738 60.05 36.703 ;
        RECT 43.076 36.666 60.004 36.749 ;
        RECT 48.596 31.146 65.525 31.228 ;
        RECT 59.958 19.784 60.004 36.749 ;
        RECT 43.03 36.712 59.958 36.795 ;
        RECT 48.642 31.1 65.571 31.182 ;
        RECT 59.912 19.83 59.958 36.795 ;
        RECT 42.984 36.758 59.912 36.841 ;
        RECT 48.688 31.054 65.617 31.136 ;
        RECT 59.866 19.876 59.912 36.841 ;
        RECT 42.938 36.804 59.866 36.887 ;
        RECT 48.734 31.008 65.663 31.09 ;
        RECT 59.82 19.922 59.866 36.887 ;
        RECT 42.892 36.85 59.82 36.933 ;
        RECT 48.78 30.962 65.709 31.044 ;
        RECT 59.774 19.968 59.82 36.933 ;
        RECT 42.846 36.896 59.774 36.979 ;
        RECT 48.826 30.916 65.755 30.998 ;
        RECT 59.728 20.014 59.774 36.979 ;
        RECT 42.8 36.942 59.728 37.025 ;
        RECT 48.872 30.87 65.801 30.952 ;
        RECT 59.682 20.06 59.728 37.025 ;
        RECT 42.754 36.988 59.682 37.071 ;
        RECT 48.918 30.824 65.847 30.906 ;
        RECT 59.636 20.106 59.682 37.071 ;
        RECT 42.708 37.034 59.636 37.117 ;
        RECT 48.964 30.778 65.893 30.86 ;
        RECT 59.59 20.152 59.636 37.117 ;
        RECT 42.662 37.08 59.59 37.163 ;
        RECT 49.01 30.732 65.939 30.814 ;
        RECT 59.544 20.198 59.59 37.163 ;
        RECT 42.616 37.126 59.544 37.209 ;
        RECT 49.056 30.686 65.985 30.768 ;
        RECT 59.498 20.244 59.544 37.209 ;
        RECT 42.57 37.172 59.498 37.255 ;
        RECT 49.102 30.64 66.031 30.722 ;
        RECT 59.452 20.29 59.498 37.255 ;
        RECT 42.524 37.218 59.452 37.301 ;
        RECT 49.148 30.594 66.077 30.676 ;
        RECT 59.406 20.336 59.452 37.301 ;
        RECT 42.478 37.264 59.406 37.347 ;
        RECT 49.194 30.548 66.123 30.63 ;
        RECT 59.36 20.382 59.406 37.347 ;
        RECT 42.432 37.31 59.36 37.393 ;
        RECT 49.24 30.502 66.169 30.584 ;
        RECT 59.314 20.428 59.36 37.393 ;
        RECT 42.386 37.356 59.314 37.439 ;
        RECT 49.286 30.456 66.215 30.538 ;
        RECT 59.268 20.474 59.314 37.439 ;
        RECT 42.34 37.402 59.268 37.485 ;
        RECT 49.332 30.41 66.261 30.492 ;
        RECT 59.222 20.52 59.268 37.485 ;
        RECT 42.294 37.448 59.222 37.531 ;
        RECT 49.378 30.364 66.307 30.446 ;
        RECT 59.176 20.566 59.222 37.531 ;
        RECT 42.248 37.494 59.176 37.577 ;
        RECT 49.424 30.318 66.353 30.4 ;
        RECT 59.13 20.612 59.176 37.577 ;
        RECT 42.202 37.54 59.13 37.623 ;
        RECT 49.47 30.272 66.399 30.354 ;
        RECT 59.084 20.658 59.13 37.623 ;
        RECT 42.156 37.586 59.084 37.669 ;
        RECT 49.516 30.226 66.445 30.308 ;
        RECT 59.038 20.704 59.084 37.669 ;
        RECT 42.11 37.632 59.038 37.715 ;
        RECT 49.562 30.18 66.491 30.262 ;
        RECT 58.992 20.75 59.038 37.715 ;
        RECT 42.064 37.678 58.992 37.761 ;
        RECT 49.608 30.134 66.537 30.216 ;
        RECT 58.946 20.796 58.992 37.761 ;
        RECT 42.018 37.724 58.946 37.807 ;
        RECT 49.654 30.088 66.583 30.17 ;
        RECT 58.9 20.842 58.946 37.807 ;
        RECT 41.972 37.77 58.9 37.853 ;
        RECT 49.7 30.042 66.629 30.124 ;
        RECT 58.854 20.888 58.9 37.853 ;
        RECT 41.926 37.816 58.854 37.899 ;
        RECT 49.746 29.996 66.675 30.078 ;
        RECT 58.808 20.934 58.854 37.899 ;
        RECT 41.88 37.862 58.808 37.945 ;
        RECT 49.792 29.95 66.721 30.032 ;
        RECT 58.762 20.98 58.808 37.945 ;
        RECT 41.834 37.908 58.762 37.991 ;
        RECT 49.838 29.904 66.767 29.986 ;
        RECT 58.716 21.026 58.762 37.991 ;
        RECT 41.788 37.954 58.716 38.037 ;
        RECT 49.884 29.858 66.813 29.94 ;
        RECT 58.67 21.072 58.716 38.037 ;
        RECT 41.742 38 58.67 38.083 ;
        RECT 49.93 29.812 66.859 29.894 ;
        RECT 58.624 21.118 58.67 38.083 ;
        RECT 41.696 38.046 58.624 38.129 ;
        RECT 49.976 29.766 66.905 29.848 ;
        RECT 58.578 21.164 58.624 38.129 ;
        RECT 41.65 38.092 58.578 38.175 ;
        RECT 50.022 29.72 66.951 29.802 ;
        RECT 58.532 21.21 58.578 38.175 ;
        RECT 41.604 38.138 58.532 38.221 ;
        RECT 50.068 29.674 66.997 29.756 ;
        RECT 58.486 21.256 58.532 38.221 ;
        RECT 41.558 38.184 58.486 38.267 ;
        RECT 50.114 29.628 67.043 29.71 ;
        RECT 58.44 21.302 58.486 38.267 ;
        RECT 41.512 38.23 58.44 38.313 ;
        RECT 50.16 29.582 67.089 29.664 ;
        RECT 58.394 21.348 58.44 38.313 ;
        RECT 41.466 38.276 58.394 38.359 ;
        RECT 50.206 29.536 67.135 29.618 ;
        RECT 58.348 21.394 58.394 38.359 ;
        RECT 41.42 38.322 58.348 38.405 ;
        RECT 50.252 29.49 67.181 29.572 ;
        RECT 58.302 21.44 58.348 38.405 ;
        RECT 41.374 38.368 58.302 38.451 ;
        RECT 50.298 29.444 67.227 29.526 ;
        RECT 58.256 21.486 58.302 38.451 ;
        RECT 41.328 38.414 58.256 38.497 ;
        RECT 50.344 29.398 67.273 29.48 ;
        RECT 58.21 21.532 58.256 38.497 ;
        RECT 41.282 38.46 58.21 38.543 ;
        RECT 50.39 29.352 67.319 29.434 ;
        RECT 58.164 21.578 58.21 38.543 ;
        RECT 41.236 38.506 58.164 38.589 ;
        RECT 50.436 29.306 67.365 29.388 ;
        RECT 58.118 21.624 58.164 38.589 ;
        RECT 41.19 38.552 58.118 38.635 ;
        RECT 50.482 29.26 67.411 29.342 ;
        RECT 58.072 21.67 58.118 38.635 ;
        RECT 41.144 38.598 58.072 38.681 ;
        RECT 50.528 29.214 67.457 29.296 ;
        RECT 58.026 21.716 58.072 38.681 ;
        RECT 41.098 38.644 58.026 38.727 ;
        RECT 50.574 29.168 67.503 29.25 ;
        RECT 57.98 21.762 58.026 38.727 ;
        RECT 41.052 38.69 57.98 38.773 ;
        RECT 50.62 29.122 67.549 29.204 ;
        RECT 57.934 21.808 57.98 38.773 ;
        RECT 41.006 38.736 57.934 38.819 ;
        RECT 50.666 29.076 67.595 29.158 ;
        RECT 57.888 21.854 57.934 38.819 ;
        RECT 40.96 38.782 57.888 38.865 ;
        RECT 50.712 29.03 67.641 29.112 ;
        RECT 57.842 21.9 57.888 38.865 ;
        RECT 40.914 38.828 57.842 38.911 ;
        RECT 50.758 28.984 67.687 29.066 ;
        RECT 57.796 21.946 57.842 38.911 ;
        RECT 40.868 38.874 57.796 38.957 ;
        RECT 50.804 28.938 110 29 ;
        RECT 57.75 21.992 57.796 38.957 ;
        RECT 40.822 38.92 57.75 39.003 ;
        RECT 50.85 28.892 110 29 ;
        RECT 57.704 22.038 57.75 39.003 ;
        RECT 40.776 38.966 57.704 39.049 ;
        RECT 50.896 28.846 110 29 ;
        RECT 57.658 22.084 57.704 39.049 ;
        RECT 40.73 39.012 57.658 39.095 ;
        RECT 50.942 28.8 110 29 ;
        RECT 57.612 22.13 57.658 39.095 ;
        RECT 40.684 39.058 57.612 39.141 ;
        RECT 50.988 28.754 110 29 ;
        RECT 57.566 22.176 57.612 39.141 ;
        RECT 40.638 39.104 57.566 39.187 ;
        RECT 51.034 28.708 110 29 ;
        RECT 57.52 22.222 57.566 39.187 ;
        RECT 40.592 39.15 57.52 39.233 ;
        RECT 51.08 28.662 110 29 ;
        RECT 57.474 22.268 57.52 39.233 ;
        RECT 40.546 39.196 57.474 39.279 ;
        RECT 51.126 28.616 110 29 ;
        RECT 57.428 22.314 57.474 39.279 ;
        RECT 40.5 39.242 57.428 39.325 ;
        RECT 51.172 28.57 110 29 ;
        RECT 57.382 22.36 57.428 39.325 ;
        RECT 40.454 39.288 57.382 39.371 ;
        RECT 51.218 28.524 110 29 ;
        RECT 57.336 22.406 57.382 39.371 ;
        RECT 40.408 39.334 57.336 39.417 ;
        RECT 51.264 28.478 110 29 ;
        RECT 57.29 22.452 57.336 39.417 ;
        RECT 40.362 39.38 57.29 39.463 ;
        RECT 51.31 28.432 110 29 ;
        RECT 57.244 22.498 57.29 39.463 ;
        RECT 40.316 39.426 57.244 39.509 ;
        RECT 51.356 28.386 110 29 ;
        RECT 57.198 22.544 57.244 39.509 ;
        RECT 40.27 39.472 57.198 39.555 ;
        RECT 51.402 28.34 110 29 ;
        RECT 57.152 22.59 57.198 39.555 ;
        RECT 40.224 39.518 57.152 39.601 ;
        RECT 51.448 28.294 110 29 ;
        RECT 57.106 22.636 57.152 39.601 ;
        RECT 40.178 39.564 57.106 39.647 ;
        RECT 51.494 28.248 110 29 ;
        RECT 57.06 22.682 57.106 39.647 ;
        RECT 40.132 39.61 57.06 39.693 ;
        RECT 51.54 28.202 110 29 ;
        RECT 57.014 22.728 57.06 39.693 ;
        RECT 40.086 39.656 57.014 39.739 ;
        RECT 51.586 28.156 110 29 ;
        RECT 56.968 22.774 57.014 39.739 ;
        RECT 40.04 39.702 56.968 39.785 ;
        RECT 51.632 28.11 110 29 ;
        RECT 56.922 22.82 56.968 39.785 ;
        RECT 39.994 39.748 56.922 39.831 ;
        RECT 51.678 28.064 110 29 ;
        RECT 56.876 22.866 56.922 39.831 ;
        RECT 39.948 39.794 56.876 39.877 ;
        RECT 51.724 28.018 110 29 ;
        RECT 56.83 22.912 56.876 39.877 ;
        RECT 39.902 39.84 56.83 39.923 ;
        RECT 51.77 27.972 110 29 ;
        RECT 56.784 22.958 56.83 39.923 ;
        RECT 39.856 39.886 56.784 39.969 ;
        RECT 51.816 27.926 110 29 ;
        RECT 56.738 23.004 56.784 39.969 ;
        RECT 39.81 39.932 56.738 40.015 ;
        RECT 51.862 27.88 110 29 ;
        RECT 56.692 23.05 56.738 40.015 ;
        RECT 39.764 39.978 56.692 40.061 ;
        RECT 51.908 27.834 110 29 ;
        RECT 56.646 23.096 56.692 40.061 ;
        RECT 39.718 40.024 56.646 40.107 ;
        RECT 51.954 27.788 110 29 ;
        RECT 56.6 23.142 56.646 40.107 ;
        RECT 39.672 40.07 56.6 40.153 ;
        RECT 52 27.742 110 29 ;
        RECT 56.554 23.188 56.6 40.153 ;
        RECT 39.626 40.116 56.554 40.199 ;
        RECT 52.046 27.696 110 29 ;
        RECT 56.508 23.234 56.554 40.199 ;
        RECT 39.58 40.162 56.508 40.245 ;
        RECT 52.092 27.65 110 29 ;
        RECT 56.462 23.28 56.508 40.245 ;
        RECT 39.534 40.208 56.462 40.291 ;
        RECT 52.138 27.604 110 29 ;
        RECT 56.416 23.326 56.462 40.291 ;
        RECT 39.488 40.254 56.416 40.337 ;
        RECT 52.184 27.558 110 29 ;
        RECT 56.37 23.372 56.416 40.337 ;
        RECT 39.442 40.3 56.37 40.383 ;
        RECT 52.23 27.512 110 29 ;
        RECT 56.324 23.418 56.37 40.383 ;
        RECT 39.396 40.346 56.324 40.429 ;
        RECT 52.276 27.466 110 29 ;
        RECT 56.278 23.464 56.324 40.429 ;
        RECT 39.35 40.392 56.278 40.475 ;
        RECT 52.322 27.42 110 29 ;
        RECT 56.232 23.51 56.278 40.475 ;
        RECT 39.304 40.438 56.232 40.521 ;
        RECT 52.368 27.374 110 29 ;
        RECT 56.186 23.556 56.232 40.521 ;
        RECT 39.258 40.484 56.186 40.567 ;
        RECT 52.414 27.328 110 29 ;
        RECT 56.14 23.602 56.186 40.567 ;
        RECT 39.212 40.53 56.14 40.613 ;
        RECT 52.46 27.282 110 29 ;
        RECT 56.094 23.648 56.14 40.613 ;
        RECT 39.166 40.576 56.094 40.659 ;
        RECT 52.506 27.236 110 29 ;
        RECT 56.048 23.694 56.094 40.659 ;
        RECT 39.12 40.622 56.048 40.705 ;
        RECT 52.552 27.19 110 29 ;
        RECT 56.002 23.74 56.048 40.705 ;
        RECT 39.074 40.668 56.002 40.751 ;
        RECT 52.598 27.144 110 29 ;
        RECT 55.956 23.786 56.002 40.751 ;
        RECT 39.028 40.714 55.956 40.797 ;
        RECT 52.644 27.098 110 29 ;
        RECT 55.91 23.832 55.956 40.797 ;
        RECT 38.982 40.76 55.91 40.843 ;
        RECT 52.69 27.052 110 29 ;
        RECT 55.864 23.878 55.91 40.843 ;
        RECT 38.936 40.806 55.864 40.889 ;
        RECT 52.736 27.006 110 29 ;
        RECT 55.818 23.924 55.864 40.889 ;
        RECT 38.89 40.852 55.818 40.935 ;
        RECT 52.782 26.96 110 29 ;
        RECT 55.772 23.97 55.818 40.935 ;
        RECT 38.844 40.898 55.772 40.981 ;
        RECT 52.828 26.914 110 29 ;
        RECT 55.726 24.016 55.772 40.981 ;
        RECT 38.798 40.944 55.726 41.027 ;
        RECT 52.874 26.868 110 29 ;
        RECT 55.68 24.062 55.726 41.027 ;
        RECT 38.752 40.99 55.68 41.073 ;
        RECT 52.92 26.822 110 29 ;
        RECT 55.634 24.108 55.68 41.073 ;
        RECT 38.706 41.036 55.634 41.119 ;
        RECT 52.966 26.776 110 29 ;
        RECT 55.588 24.154 55.634 41.119 ;
        RECT 38.66 41.082 55.588 41.165 ;
        RECT 53.012 26.73 110 29 ;
        RECT 55.542 24.2 55.588 41.165 ;
        RECT 38.614 41.128 55.542 41.211 ;
        RECT 53.058 26.684 110 29 ;
        RECT 55.496 24.246 55.542 41.211 ;
        RECT 38.568 41.174 55.496 41.257 ;
        RECT 53.104 26.638 110 29 ;
        RECT 55.45 24.292 55.496 41.257 ;
        RECT 38.522 41.22 55.45 41.303 ;
        RECT 53.15 26.592 110 29 ;
        RECT 55.404 24.338 55.45 41.303 ;
        RECT 38.476 41.266 55.404 41.349 ;
        RECT 53.196 26.546 110 29 ;
        RECT 55.358 24.384 55.404 41.349 ;
        RECT 38.43 41.312 55.358 41.395 ;
        RECT 53.242 26.5 110 29 ;
        RECT 55.312 24.43 55.358 41.395 ;
        RECT 38.384 41.358 55.312 41.441 ;
        RECT 53.288 26.454 110 29 ;
        RECT 55.266 24.476 55.312 41.441 ;
        RECT 38.338 41.404 55.266 41.487 ;
        RECT 53.334 26.408 110 29 ;
        RECT 55.22 24.522 55.266 41.487 ;
        RECT 38.292 41.45 55.22 41.533 ;
        RECT 53.38 26.362 110 29 ;
        RECT 55.174 24.568 55.22 41.533 ;
        RECT 38.246 41.496 55.174 41.579 ;
        RECT 53.426 26.316 110 29 ;
        RECT 55.128 24.614 55.174 41.579 ;
        RECT 38.2 41.542 55.128 41.625 ;
        RECT 53.472 26.27 110 29 ;
        RECT 55.082 24.66 55.128 41.625 ;
        RECT 38.154 41.588 55.082 41.671 ;
        RECT 53.518 26.224 110 29 ;
        RECT 55.036 24.706 55.082 41.671 ;
        RECT 38.108 41.634 55.036 41.717 ;
        RECT 53.564 26.178 110 29 ;
        RECT 54.99 24.752 55.036 41.717 ;
        RECT 38.062 41.68 54.99 41.763 ;
        RECT 53.61 26.132 110 29 ;
        RECT 54.944 24.798 54.99 41.763 ;
        RECT 38.016 41.726 54.944 41.809 ;
        RECT 53.656 26.086 110 29 ;
        RECT 54.898 24.844 54.944 41.809 ;
        RECT 37.97 41.772 54.898 41.855 ;
        RECT 53.702 26.04 110 29 ;
        RECT 54.852 24.89 54.898 41.855 ;
        RECT 37.924 41.818 54.852 41.901 ;
        RECT 53.748 25.994 110 29 ;
        RECT 54.806 24.936 54.852 41.901 ;
        RECT 37.878 41.864 54.806 41.947 ;
        RECT 53.794 25.948 110 29 ;
        RECT 54.76 24.982 54.806 41.947 ;
        RECT 37.832 41.91 54.76 41.993 ;
        RECT 53.84 25.902 110 29 ;
        RECT 54.714 25.028 54.76 41.993 ;
        RECT 37.786 41.956 54.714 42.039 ;
        RECT 53.886 25.856 110 29 ;
        RECT 54.668 25.074 54.714 42.039 ;
        RECT 37.74 42.002 54.668 42.085 ;
        RECT 53.932 25.81 110 29 ;
        RECT 54.622 25.12 54.668 42.085 ;
        RECT 37.694 42.048 54.622 42.131 ;
        RECT 53.978 25.764 110 29 ;
        RECT 54.576 25.166 54.622 42.131 ;
        RECT 37.648 42.094 54.576 42.177 ;
        RECT 54.024 25.718 110 29 ;
        RECT 54.53 25.212 54.576 42.177 ;
        RECT 37.602 42.14 54.53 42.223 ;
        RECT 54.07 25.672 110 29 ;
        RECT 54.484 25.258 54.53 42.223 ;
        RECT 37.556 42.186 54.484 42.269 ;
        RECT 54.116 25.626 110 29 ;
        RECT 54.438 25.304 54.484 42.269 ;
        RECT 37.51 42.232 54.438 42.315 ;
        RECT 54.162 25.58 110 29 ;
        RECT 54.392 25.35 54.438 42.315 ;
        RECT 37.464 42.278 54.392 42.361 ;
        RECT 54.208 25.534 110 29 ;
        RECT 54.346 25.396 54.392 42.361 ;
        RECT 37.418 42.324 54.346 42.407 ;
        RECT 54.254 25.488 110 29 ;
        RECT 54.3 25.442 54.346 42.407 ;
        RECT 37.372 42.37 54.3 42.453 ;
        RECT 37.326 42.416 54.254 42.499 ;
        RECT 37.28 42.462 54.208 42.545 ;
        RECT 37.234 42.508 54.162 42.591 ;
        RECT 37.188 42.554 54.116 42.637 ;
        RECT 37.142 42.6 54.07 42.683 ;
        RECT 37.096 42.646 54.024 42.729 ;
        RECT 37.05 42.692 53.978 42.775 ;
        RECT 37.004 42.738 53.932 42.821 ;
        RECT 36.958 42.784 53.886 42.867 ;
        RECT 36.912 42.83 53.84 42.913 ;
        RECT 36.866 42.876 53.794 42.959 ;
        RECT 36.82 42.922 53.748 43.005 ;
        RECT 36.774 42.968 53.702 43.051 ;
        RECT 36.728 43.014 53.656 43.097 ;
        RECT 36.682 43.06 53.61 43.143 ;
        RECT 36.636 43.106 53.564 43.189 ;
        RECT 36.59 43.152 53.518 43.235 ;
        RECT 36.544 43.198 53.472 43.281 ;
        RECT 36.498 43.244 53.426 43.327 ;
        RECT 36.452 43.29 53.38 43.373 ;
        RECT 36.406 43.336 53.334 43.419 ;
        RECT 36.36 43.382 53.288 43.465 ;
        RECT 36.314 43.428 53.242 43.511 ;
        RECT 36.268 43.474 53.196 43.557 ;
        RECT 36.222 43.52 53.15 43.603 ;
        RECT 36.176 43.566 53.104 43.649 ;
        RECT 36.13 43.612 53.058 43.695 ;
        RECT 36.084 43.658 53.012 43.741 ;
        RECT 36.038 43.704 52.966 43.787 ;
        RECT 35.992 43.75 52.92 43.833 ;
        RECT 35.946 43.796 52.874 43.879 ;
        RECT 35.9 43.842 52.828 43.925 ;
        RECT 35.854 43.888 52.782 43.971 ;
        RECT 35.808 43.934 52.736 44.017 ;
        RECT 35.762 43.98 52.69 44.063 ;
        RECT 35.716 44.026 52.644 44.109 ;
        RECT 35.67 44.072 52.598 44.155 ;
        RECT 35.624 44.118 52.552 44.201 ;
        RECT 35.578 44.164 52.506 44.247 ;
        RECT 35.532 44.21 52.46 44.293 ;
        RECT 35.486 44.256 52.414 44.339 ;
        RECT 35.44 44.302 52.368 44.385 ;
        RECT 35.394 44.348 52.322 44.431 ;
        RECT 35.348 44.394 52.276 44.477 ;
        RECT 35.302 44.44 52.23 44.523 ;
        RECT 35.256 44.486 52.184 44.569 ;
        RECT 35.21 44.532 52.138 44.615 ;
        RECT 35.164 44.578 52.092 44.661 ;
        RECT 35.118 44.624 52.046 44.707 ;
        RECT 35.072 44.67 52 44.753 ;
        RECT 35.026 44.716 51.954 44.799 ;
        RECT 34.98 44.762 51.908 44.845 ;
        RECT 34.934 44.808 51.862 44.891 ;
        RECT 34.888 44.854 51.816 44.937 ;
        RECT 34.842 44.9 51.77 44.983 ;
        RECT 34.796 44.946 51.724 45.029 ;
        RECT 34.75 44.992 51.678 45.075 ;
        RECT 34.704 45.038 51.632 45.121 ;
        RECT 34.658 45.084 51.586 45.167 ;
        RECT 34.612 45.13 51.54 45.213 ;
        RECT 34.566 45.176 51.494 45.259 ;
        RECT 34.52 45.222 51.448 45.305 ;
        RECT 34.474 45.268 51.402 45.351 ;
        RECT 34.428 45.314 51.356 45.397 ;
        RECT 34.382 45.36 51.31 45.443 ;
        RECT 34.336 45.406 51.264 45.489 ;
        RECT 34.29 45.452 51.218 45.535 ;
        RECT 34.244 45.498 51.172 45.581 ;
        RECT 34.198 45.544 51.126 45.627 ;
        RECT 34.152 45.59 51.08 45.673 ;
        RECT 34.106 45.636 51.034 45.719 ;
        RECT 34.06 45.682 50.988 45.765 ;
        RECT 34.014 45.728 50.942 45.811 ;
        RECT 33.968 45.774 50.896 45.857 ;
        RECT 33.922 45.82 50.85 45.903 ;
        RECT 33.876 45.866 50.804 45.949 ;
        RECT 33.83 45.912 50.758 45.995 ;
        RECT 33.784 45.958 50.712 46.041 ;
        RECT 33.738 46.004 50.666 46.087 ;
        RECT 33.692 46.05 50.62 46.133 ;
        RECT 33.646 46.096 50.574 46.179 ;
        RECT 33.6 46.142 50.528 46.225 ;
        RECT 33.554 46.188 50.482 46.271 ;
        RECT 33.508 46.234 50.436 46.317 ;
        RECT 33.462 46.28 50.39 46.363 ;
        RECT 33.416 46.326 50.344 46.409 ;
        RECT 33.37 46.372 50.298 46.455 ;
        RECT 33.324 46.418 50.252 46.501 ;
        RECT 33.278 46.464 50.206 46.547 ;
        RECT 33.232 46.51 50.16 46.593 ;
        RECT 33.186 46.556 50.114 46.639 ;
        RECT 33.14 46.602 50.068 46.685 ;
        RECT 33.094 46.648 50.022 46.731 ;
        RECT 33.048 46.694 49.976 46.777 ;
        RECT 33.002 46.74 49.93 46.823 ;
        RECT 32.956 46.786 49.884 46.869 ;
        RECT 32.91 46.832 49.838 46.915 ;
        RECT 32.864 46.878 49.792 46.961 ;
        RECT 32.818 46.924 49.746 47.007 ;
        RECT 32.772 46.97 49.7 47.053 ;
        RECT 32.726 47.016 49.654 47.099 ;
        RECT 32.68 47.062 49.608 47.145 ;
        RECT 32.634 47.108 49.562 47.191 ;
        RECT 32.588 47.154 49.516 47.237 ;
        RECT 32.542 47.2 49.47 47.283 ;
        RECT 32.496 47.246 49.424 47.329 ;
        RECT 32.45 47.292 49.378 47.375 ;
        RECT 32.404 47.338 49.332 47.421 ;
        RECT 32.358 47.384 49.286 47.467 ;
        RECT 32.312 47.43 49.24 47.513 ;
        RECT 32.266 47.476 49.194 47.559 ;
        RECT 32.22 47.522 49.148 47.605 ;
        RECT 32.174 47.568 49.102 47.651 ;
        RECT 32.128 47.614 49.056 47.697 ;
        RECT 32.082 47.66 49.01 47.743 ;
        RECT 32.036 47.706 48.964 47.789 ;
        RECT 31.99 47.752 48.918 47.835 ;
        RECT 31.944 47.798 48.872 47.881 ;
        RECT 31.898 47.844 48.826 47.927 ;
        RECT 31.852 47.89 48.78 47.973 ;
        RECT 31.806 47.936 48.734 48.019 ;
        RECT 31.76 47.982 48.688 48.065 ;
        RECT 31.714 48.028 48.642 48.111 ;
        RECT 31.668 48.074 48.596 48.157 ;
        RECT 31.622 48.12 48.55 48.203 ;
        RECT 31.576 48.166 48.504 48.249 ;
        RECT 31.53 48.212 48.458 48.295 ;
        RECT 31.484 48.258 48.412 48.341 ;
        RECT 31.438 48.304 48.366 48.387 ;
        RECT 31.392 48.35 48.32 48.433 ;
        RECT 31.346 48.396 48.274 48.479 ;
        RECT 31.3 48.442 48.228 48.525 ;
        RECT 31.254 48.488 48.182 48.571 ;
        RECT 31.208 48.534 48.136 48.617 ;
        RECT 31.162 48.58 48.09 48.663 ;
        RECT 31.116 48.626 48.044 48.709 ;
        RECT 31.07 48.672 47.998 48.755 ;
        RECT 31.024 48.718 47.952 48.801 ;
        RECT 30.978 48.764 47.906 48.847 ;
        RECT 30.932 48.81 47.86 48.893 ;
        RECT 30.886 48.856 47.814 48.939 ;
        RECT 30.84 48.902 47.768 48.985 ;
        RECT 30.794 48.948 47.722 49.031 ;
        RECT 30.748 48.994 47.676 49.077 ;
        RECT 30.702 49.04 47.63 49.123 ;
        RECT 30.656 49.086 47.584 49.169 ;
        RECT 30.61 49.132 47.538 49.215 ;
        RECT 30.564 49.178 47.492 49.261 ;
        RECT 30.518 49.224 47.446 49.307 ;
        RECT 30.472 49.27 47.4 49.353 ;
        RECT 30.426 49.316 47.354 49.399 ;
        RECT 30.38 49.362 47.308 49.445 ;
        RECT 30.334 49.408 47.262 49.491 ;
        RECT 30.288 49.454 47.216 49.537 ;
        RECT 30.242 49.5 47.17 49.583 ;
        RECT 30.196 49.546 47.124 49.629 ;
        RECT 30.15 49.592 47.078 49.675 ;
        RECT 30.104 49.638 47.032 49.721 ;
        RECT 30.058 49.684 46.986 49.767 ;
        RECT 30.012 49.73 46.94 49.813 ;
        RECT 29.966 49.776 46.894 49.859 ;
        RECT 29.92 49.822 46.848 49.905 ;
        RECT 29.874 49.868 46.802 49.951 ;
        RECT 29.828 49.914 46.756 49.997 ;
        RECT 29.782 49.96 46.71 50.043 ;
        RECT 29.736 50.006 46.664 50.089 ;
        RECT 29.69 50.052 46.618 50.135 ;
        RECT 29.644 50.098 46.572 50.181 ;
        RECT 29.598 50.144 46.526 50.227 ;
        RECT 29.552 50.19 46.48 50.273 ;
        RECT 29.506 50.236 46.434 50.319 ;
        RECT 29.46 50.282 46.388 50.365 ;
        RECT 29.414 50.328 46.342 50.411 ;
        RECT 29.368 50.374 46.296 50.457 ;
        RECT 29.322 50.42 46.25 50.503 ;
        RECT 29.276 50.466 46.204 50.549 ;
        RECT 29.23 50.512 46.158 50.595 ;
        RECT 29.184 50.558 46.112 50.641 ;
        RECT 29.138 50.604 46.066 50.687 ;
        RECT 29.092 50.65 46.02 50.733 ;
        RECT 29.046 50.696 45.974 50.779 ;
        RECT 29 50.742 45.928 50.825 ;
        RECT 28.96 50.785 45.882 50.871 ;
        RECT 28.914 50.828 45.836 50.917 ;
        RECT 28.868 50.874 45.79 50.963 ;
        RECT 28.822 50.92 45.744 51.009 ;
        RECT 28.776 50.966 45.698 51.055 ;
        RECT 28.73 51.012 45.652 51.101 ;
        RECT 28.684 51.058 45.606 51.147 ;
        RECT 28.638 51.104 45.56 51.193 ;
        RECT 28.592 51.15 45.514 51.239 ;
        RECT 28.546 51.196 45.468 51.285 ;
        RECT 28.5 51.242 45.422 51.331 ;
        RECT 28.454 51.288 45.376 51.377 ;
        RECT 28.408 51.334 45.33 51.423 ;
        RECT 28.362 51.38 45.284 51.469 ;
        RECT 56.015 3.5 110 15.5 ;
        RECT 39.098 20.394 56.061 20.442 ;
        RECT 55.98 3.517 56.015 20.483 ;
        RECT 39.052 20.44 55.98 20.523 ;
        RECT 39.144 20.348 56.107 20.396 ;
        RECT 55.934 3.558 55.98 20.523 ;
        RECT 39.006 20.486 55.934 20.569 ;
        RECT 39.19 20.302 56.153 20.35 ;
        RECT 55.888 3.604 55.934 20.569 ;
        RECT 38.96 20.532 55.888 20.615 ;
        RECT 39.236 20.256 56.199 20.304 ;
        RECT 55.842 3.65 55.888 20.615 ;
        RECT 38.914 20.578 55.842 20.661 ;
        RECT 39.282 20.21 56.245 20.258 ;
        RECT 55.796 3.696 55.842 20.661 ;
        RECT 38.868 20.624 55.796 20.707 ;
        RECT 39.328 20.164 56.291 20.212 ;
        RECT 55.75 3.742 55.796 20.707 ;
        RECT 38.822 20.67 55.75 20.753 ;
        RECT 39.374 20.118 56.337 20.166 ;
        RECT 55.704 3.788 55.75 20.753 ;
        RECT 38.776 20.716 55.704 20.799 ;
        RECT 39.42 20.072 56.383 20.12 ;
        RECT 55.658 3.834 55.704 20.799 ;
        RECT 38.73 20.762 55.658 20.845 ;
        RECT 39.466 20.026 56.429 20.074 ;
        RECT 55.612 3.88 55.658 20.845 ;
        RECT 38.684 20.808 55.612 20.891 ;
        RECT 39.512 19.98 56.475 20.028 ;
        RECT 55.566 3.926 55.612 20.891 ;
        RECT 38.638 20.854 55.566 20.937 ;
        RECT 39.558 19.934 56.521 19.982 ;
        RECT 55.52 3.972 55.566 20.937 ;
        RECT 38.592 20.9 55.52 20.983 ;
        RECT 39.604 19.888 56.567 19.936 ;
        RECT 55.474 4.018 55.52 20.983 ;
        RECT 38.546 20.946 55.474 21.029 ;
        RECT 39.65 19.842 56.613 19.89 ;
        RECT 55.428 4.064 55.474 21.029 ;
        RECT 38.5 20.992 55.428 21.075 ;
        RECT 39.696 19.796 56.659 19.844 ;
        RECT 55.382 4.11 55.428 21.075 ;
        RECT 38.454 21.038 55.382 21.121 ;
        RECT 39.742 19.75 56.705 19.798 ;
        RECT 55.336 4.156 55.382 21.121 ;
        RECT 38.408 21.084 55.336 21.167 ;
        RECT 39.788 19.704 56.751 19.752 ;
        RECT 55.29 4.202 55.336 21.167 ;
        RECT 38.362 21.13 55.29 21.213 ;
        RECT 39.834 19.658 56.797 19.706 ;
        RECT 55.244 4.248 55.29 21.213 ;
        RECT 38.316 21.176 55.244 21.259 ;
        RECT 39.88 19.612 56.843 19.66 ;
        RECT 55.198 4.294 55.244 21.259 ;
        RECT 38.27 21.222 55.198 21.305 ;
        RECT 39.926 19.566 56.889 19.614 ;
        RECT 55.152 4.34 55.198 21.305 ;
        RECT 38.224 21.268 55.152 21.351 ;
        RECT 39.972 19.52 56.935 19.568 ;
        RECT 55.106 4.386 55.152 21.351 ;
        RECT 38.178 21.314 55.106 21.397 ;
        RECT 40.018 19.474 56.981 19.522 ;
        RECT 55.06 4.432 55.106 21.397 ;
        RECT 38.132 21.36 55.06 21.443 ;
        RECT 40.064 19.428 57.027 19.476 ;
        RECT 55.014 4.478 55.06 21.443 ;
        RECT 38.086 21.406 55.014 21.489 ;
        RECT 40.11 19.382 57.073 19.43 ;
        RECT 54.968 4.524 55.014 21.489 ;
        RECT 38.04 21.452 54.968 21.535 ;
        RECT 40.156 19.336 57.119 19.384 ;
        RECT 54.922 4.57 54.968 21.535 ;
        RECT 37.994 21.498 54.922 21.581 ;
        RECT 40.202 19.29 57.165 19.338 ;
        RECT 54.876 4.616 54.922 21.581 ;
        RECT 37.948 21.544 54.876 21.627 ;
        RECT 40.248 19.244 57.211 19.292 ;
        RECT 54.83 4.662 54.876 21.627 ;
        RECT 37.902 21.59 54.83 21.673 ;
        RECT 40.294 19.198 57.257 19.246 ;
        RECT 54.784 4.708 54.83 21.673 ;
        RECT 37.856 21.636 54.784 21.719 ;
        RECT 40.34 19.152 57.303 19.2 ;
        RECT 54.738 4.754 54.784 21.719 ;
        RECT 37.81 21.682 54.738 21.765 ;
        RECT 40.386 19.106 57.349 19.154 ;
        RECT 54.692 4.8 54.738 21.765 ;
        RECT 37.764 21.728 54.692 21.811 ;
        RECT 40.432 19.06 57.395 19.108 ;
        RECT 54.646 4.846 54.692 21.811 ;
        RECT 37.718 21.774 54.646 21.857 ;
        RECT 40.478 19.014 57.441 19.062 ;
        RECT 54.6 4.892 54.646 21.857 ;
        RECT 37.672 21.82 54.6 21.903 ;
        RECT 40.524 18.968 57.487 19.016 ;
        RECT 54.554 4.938 54.6 21.903 ;
        RECT 37.626 21.866 54.554 21.949 ;
        RECT 40.57 18.922 57.533 18.97 ;
        RECT 54.508 4.984 54.554 21.949 ;
        RECT 37.58 21.912 54.508 21.995 ;
        RECT 40.616 18.876 57.579 18.924 ;
        RECT 54.462 5.03 54.508 21.995 ;
        RECT 37.534 21.958 54.462 22.041 ;
        RECT 40.662 18.83 57.625 18.878 ;
        RECT 54.416 5.076 54.462 22.041 ;
        RECT 37.488 22.004 54.416 22.087 ;
        RECT 40.708 18.784 57.671 18.832 ;
        RECT 54.37 5.122 54.416 22.087 ;
        RECT 37.442 22.05 54.37 22.133 ;
        RECT 40.754 18.738 57.717 18.786 ;
        RECT 54.324 5.168 54.37 22.133 ;
        RECT 37.396 22.096 54.324 22.179 ;
        RECT 40.8 18.692 57.763 18.74 ;
        RECT 54.278 5.214 54.324 22.179 ;
        RECT 37.35 22.142 54.278 22.225 ;
        RECT 40.846 18.646 57.809 18.694 ;
        RECT 54.232 5.26 54.278 22.225 ;
        RECT 37.304 22.188 54.232 22.271 ;
        RECT 40.892 18.6 57.855 18.648 ;
        RECT 54.186 5.306 54.232 22.271 ;
        RECT 37.258 22.234 54.186 22.317 ;
        RECT 40.938 18.554 57.901 18.602 ;
        RECT 54.14 5.352 54.186 22.317 ;
        RECT 37.212 22.28 54.14 22.363 ;
        RECT 40.984 18.508 57.947 18.556 ;
        RECT 54.094 5.398 54.14 22.363 ;
        RECT 37.166 22.326 54.094 22.409 ;
        RECT 41.03 18.462 57.993 18.51 ;
        RECT 54.048 5.444 54.094 22.409 ;
        RECT 37.12 22.372 54.048 22.455 ;
        RECT 41.076 18.416 58.039 18.464 ;
        RECT 54.002 5.49 54.048 22.455 ;
        RECT 37.074 22.418 54.002 22.501 ;
        RECT 41.122 18.37 58.085 18.418 ;
        RECT 53.956 5.536 54.002 22.501 ;
        RECT 37.028 22.464 53.956 22.547 ;
        RECT 41.168 18.324 58.131 18.372 ;
        RECT 53.91 5.582 53.956 22.547 ;
        RECT 36.982 22.51 53.91 22.593 ;
        RECT 41.214 18.278 58.177 18.326 ;
        RECT 53.864 5.628 53.91 22.593 ;
        RECT 36.936 22.556 53.864 22.639 ;
        RECT 41.26 18.232 58.223 18.28 ;
        RECT 53.818 5.674 53.864 22.639 ;
        RECT 36.89 22.602 53.818 22.685 ;
        RECT 41.306 18.186 58.269 18.234 ;
        RECT 53.772 5.72 53.818 22.685 ;
        RECT 36.844 22.648 53.772 22.731 ;
        RECT 41.352 18.14 58.315 18.188 ;
        RECT 53.726 5.766 53.772 22.731 ;
        RECT 36.798 22.694 53.726 22.777 ;
        RECT 41.398 18.094 58.361 18.142 ;
        RECT 53.68 5.812 53.726 22.777 ;
        RECT 36.752 22.74 53.68 22.823 ;
        RECT 41.444 18.048 58.407 18.096 ;
        RECT 53.634 5.858 53.68 22.823 ;
        RECT 36.706 22.786 53.634 22.869 ;
        RECT 41.49 18.002 58.453 18.05 ;
        RECT 53.588 5.904 53.634 22.869 ;
        RECT 36.66 22.832 53.588 22.915 ;
        RECT 41.536 17.956 58.499 18.004 ;
        RECT 53.542 5.95 53.588 22.915 ;
        RECT 36.614 22.878 53.542 22.961 ;
        RECT 41.582 17.91 58.545 17.958 ;
        RECT 53.496 5.996 53.542 22.961 ;
        RECT 36.568 22.924 53.496 23.007 ;
        RECT 41.628 17.864 58.591 17.912 ;
        RECT 53.45 6.042 53.496 23.007 ;
        RECT 36.522 22.97 53.45 23.053 ;
        RECT 41.674 17.818 58.637 17.866 ;
        RECT 53.404 6.088 53.45 23.053 ;
        RECT 36.476 23.016 53.404 23.099 ;
        RECT 41.72 17.772 58.683 17.82 ;
        RECT 53.358 6.134 53.404 23.099 ;
        RECT 36.43 23.062 53.358 23.145 ;
        RECT 41.766 17.726 58.729 17.774 ;
        RECT 53.312 6.18 53.358 23.145 ;
        RECT 36.384 23.108 53.312 23.191 ;
        RECT 41.812 17.68 58.775 17.728 ;
        RECT 53.266 6.226 53.312 23.191 ;
        RECT 36.338 23.154 53.266 23.237 ;
        RECT 41.858 17.634 58.821 17.682 ;
        RECT 53.22 6.272 53.266 23.237 ;
        RECT 36.292 23.2 53.22 23.283 ;
        RECT 41.904 17.588 58.867 17.636 ;
        RECT 53.174 6.318 53.22 23.283 ;
        RECT 36.246 23.246 53.174 23.329 ;
        RECT 41.95 17.542 58.913 17.59 ;
        RECT 53.128 6.364 53.174 23.329 ;
        RECT 36.2 23.292 53.128 23.375 ;
        RECT 41.996 17.496 58.959 17.544 ;
        RECT 53.082 6.41 53.128 23.375 ;
        RECT 36.154 23.338 53.082 23.421 ;
        RECT 42.042 17.45 59.005 17.498 ;
        RECT 53.036 6.456 53.082 23.421 ;
        RECT 36.108 23.384 53.036 23.467 ;
        RECT 42.088 17.404 59.051 17.452 ;
        RECT 52.99 6.502 53.036 23.467 ;
        RECT 36.062 23.43 52.99 23.513 ;
        RECT 42.134 17.358 59.097 17.406 ;
        RECT 52.944 6.548 52.99 23.513 ;
        RECT 36.016 23.476 52.944 23.559 ;
        RECT 42.18 17.312 59.143 17.36 ;
        RECT 52.898 6.594 52.944 23.559 ;
        RECT 35.97 23.522 52.898 23.605 ;
        RECT 42.226 17.266 59.189 17.314 ;
        RECT 52.852 6.64 52.898 23.605 ;
        RECT 35.924 23.568 52.852 23.651 ;
        RECT 42.272 17.22 59.235 17.268 ;
        RECT 52.806 6.686 52.852 23.651 ;
        RECT 35.878 23.614 52.806 23.697 ;
        RECT 42.318 17.174 59.281 17.222 ;
        RECT 52.76 6.732 52.806 23.697 ;
        RECT 35.832 23.66 52.76 23.743 ;
        RECT 42.364 17.128 59.327 17.176 ;
        RECT 52.714 6.778 52.76 23.743 ;
        RECT 35.786 23.706 52.714 23.789 ;
        RECT 42.41 17.082 59.373 17.13 ;
        RECT 52.668 6.824 52.714 23.789 ;
        RECT 35.74 23.752 52.668 23.835 ;
        RECT 42.456 17.036 59.419 17.084 ;
        RECT 52.622 6.87 52.668 23.835 ;
        RECT 35.694 23.798 52.622 23.881 ;
        RECT 42.502 16.99 59.465 17.038 ;
        RECT 52.576 6.916 52.622 23.881 ;
        RECT 35.648 23.844 52.576 23.927 ;
        RECT 42.548 16.944 59.511 16.992 ;
        RECT 52.53 6.962 52.576 23.927 ;
        RECT 35.602 23.89 52.53 23.973 ;
        RECT 42.594 16.898 59.557 16.946 ;
        RECT 52.484 7.008 52.53 23.973 ;
        RECT 35.556 23.936 52.484 24.019 ;
        RECT 42.64 16.852 59.603 16.9 ;
        RECT 52.438 7.054 52.484 24.019 ;
        RECT 35.51 23.982 52.438 24.065 ;
        RECT 42.686 16.806 59.649 16.854 ;
        RECT 52.392 7.1 52.438 24.065 ;
        RECT 35.464 24.028 52.392 24.111 ;
        RECT 42.732 16.76 59.695 16.808 ;
        RECT 52.346 7.146 52.392 24.111 ;
        RECT 35.418 24.074 52.346 24.157 ;
        RECT 42.778 16.714 59.741 16.762 ;
        RECT 52.3 7.192 52.346 24.157 ;
        RECT 35.372 24.12 52.3 24.203 ;
        RECT 42.824 16.668 59.787 16.716 ;
        RECT 52.254 7.238 52.3 24.203 ;
        RECT 35.326 24.166 52.254 24.249 ;
        RECT 42.87 16.622 59.833 16.67 ;
        RECT 52.208 7.284 52.254 24.249 ;
        RECT 35.28 24.212 52.208 24.295 ;
        RECT 42.916 16.576 59.879 16.624 ;
        RECT 52.162 7.33 52.208 24.295 ;
        RECT 35.234 24.258 52.162 24.341 ;
        RECT 42.962 16.53 59.925 16.578 ;
        RECT 52.116 7.376 52.162 24.341 ;
        RECT 35.188 24.304 52.116 24.387 ;
        RECT 43.008 16.484 59.971 16.532 ;
        RECT 52.07 7.422 52.116 24.387 ;
        RECT 35.142 24.35 52.07 24.433 ;
        RECT 43.054 16.438 60.017 16.486 ;
        RECT 52.024 7.468 52.07 24.433 ;
        RECT 35.096 24.396 52.024 24.479 ;
        RECT 43.1 16.392 60.063 16.44 ;
        RECT 51.978 7.514 52.024 24.479 ;
        RECT 35.05 24.442 51.978 24.525 ;
        RECT 43.146 16.346 60.109 16.394 ;
        RECT 51.932 7.56 51.978 24.525 ;
        RECT 35.004 24.488 51.932 24.571 ;
        RECT 43.192 16.3 60.155 16.348 ;
        RECT 51.886 7.606 51.932 24.571 ;
        RECT 34.958 24.534 51.886 24.617 ;
        RECT 43.238 16.254 60.201 16.302 ;
        RECT 51.84 7.652 51.886 24.617 ;
        RECT 34.912 24.58 51.84 24.663 ;
        RECT 43.284 16.208 60.247 16.256 ;
        RECT 51.794 7.698 51.84 24.663 ;
        RECT 34.866 24.626 51.794 24.709 ;
        RECT 43.33 16.162 60.293 16.21 ;
        RECT 51.748 7.744 51.794 24.709 ;
        RECT 34.82 24.672 51.748 24.755 ;
        RECT 43.376 16.116 60.339 16.164 ;
        RECT 51.702 7.79 51.748 24.755 ;
        RECT 34.774 24.718 51.702 24.801 ;
        RECT 43.422 16.07 60.385 16.118 ;
        RECT 51.656 7.836 51.702 24.801 ;
        RECT 34.728 24.764 51.656 24.847 ;
        RECT 43.468 16.024 60.431 16.072 ;
        RECT 51.61 7.882 51.656 24.847 ;
        RECT 34.682 24.81 51.61 24.893 ;
        RECT 43.514 15.978 60.477 16.026 ;
        RECT 51.564 7.928 51.61 24.893 ;
        RECT 34.636 24.856 51.564 24.939 ;
        RECT 43.56 15.932 60.523 15.98 ;
        RECT 51.518 7.974 51.564 24.939 ;
        RECT 34.59 24.902 51.518 24.985 ;
        RECT 43.606 15.886 60.569 15.934 ;
        RECT 51.472 8.02 51.518 24.985 ;
        RECT 34.544 24.948 51.472 25.031 ;
        RECT 43.652 15.84 60.615 15.888 ;
        RECT 51.426 8.066 51.472 25.031 ;
        RECT 34.498 24.994 51.426 25.077 ;
        RECT 43.698 15.794 60.661 15.842 ;
        RECT 51.38 8.112 51.426 25.077 ;
        RECT 34.452 25.04 51.38 25.123 ;
        RECT 43.744 15.748 60.707 15.796 ;
        RECT 51.334 8.158 51.38 25.123 ;
        RECT 34.406 25.086 51.334 25.169 ;
        RECT 43.79 15.702 60.753 15.75 ;
        RECT 51.288 8.204 51.334 25.169 ;
        RECT 34.36 25.132 51.288 25.215 ;
        RECT 43.836 15.656 60.799 15.704 ;
        RECT 51.242 8.25 51.288 25.215 ;
        RECT 34.314 25.178 51.242 25.261 ;
        RECT 43.882 15.61 60.845 15.658 ;
        RECT 51.196 8.296 51.242 25.261 ;
        RECT 34.268 25.224 51.196 25.307 ;
        RECT 43.928 15.564 60.891 15.612 ;
        RECT 51.15 8.342 51.196 25.307 ;
        RECT 34.222 25.27 51.15 25.353 ;
        RECT 43.974 15.518 60.937 15.566 ;
        RECT 51.104 8.388 51.15 25.353 ;
        RECT 34.176 25.316 51.104 25.399 ;
        RECT 44.02 15.472 60.98 15.522 ;
        RECT 51.058 8.434 51.104 25.399 ;
        RECT 34.13 25.362 51.058 25.445 ;
        RECT 44.066 15.426 110 15.5 ;
        RECT 51.012 8.48 51.058 25.445 ;
        RECT 34.084 25.408 51.012 25.491 ;
        RECT 44.112 15.38 110 15.5 ;
        RECT 50.966 8.526 51.012 25.491 ;
        RECT 34.038 25.454 50.966 25.537 ;
        RECT 44.158 15.334 110 15.5 ;
        RECT 50.92 8.572 50.966 25.537 ;
        RECT 33.992 25.5 50.92 25.583 ;
        RECT 44.204 15.288 110 15.5 ;
        RECT 50.874 8.618 50.92 25.583 ;
        RECT 33.946 25.546 50.874 25.629 ;
        RECT 44.25 15.242 110 15.5 ;
        RECT 50.828 8.664 50.874 25.629 ;
        RECT 33.9 25.592 50.828 25.675 ;
        RECT 44.296 15.196 110 15.5 ;
        RECT 50.782 8.71 50.828 25.675 ;
        RECT 33.854 25.638 50.782 25.721 ;
        RECT 44.342 15.15 110 15.5 ;
        RECT 50.736 8.756 50.782 25.721 ;
        RECT 33.808 25.684 50.736 25.767 ;
        RECT 44.388 15.104 110 15.5 ;
        RECT 50.69 8.802 50.736 25.767 ;
        RECT 33.762 25.73 50.69 25.813 ;
        RECT 44.434 15.058 110 15.5 ;
        RECT 50.644 8.848 50.69 25.813 ;
        RECT 33.716 25.776 50.644 25.859 ;
        RECT 44.48 15.012 110 15.5 ;
        RECT 50.598 8.894 50.644 25.859 ;
        RECT 33.67 25.822 50.598 25.905 ;
        RECT 44.526 14.966 110 15.5 ;
        RECT 50.552 8.94 50.598 25.905 ;
        RECT 33.624 25.868 50.552 25.951 ;
        RECT 44.572 14.92 110 15.5 ;
        RECT 50.506 8.986 50.552 25.951 ;
        RECT 33.578 25.914 50.506 25.997 ;
        RECT 44.618 14.874 110 15.5 ;
        RECT 50.46 9.032 50.506 25.997 ;
        RECT 33.532 25.96 50.46 26.043 ;
        RECT 44.664 14.828 110 15.5 ;
        RECT 50.414 9.078 50.46 26.043 ;
        RECT 33.486 26.006 50.414 26.089 ;
        RECT 44.71 14.782 110 15.5 ;
        RECT 50.368 9.124 50.414 26.089 ;
        RECT 33.44 26.052 50.368 26.135 ;
        RECT 44.756 14.736 110 15.5 ;
        RECT 50.322 9.17 50.368 26.135 ;
        RECT 33.394 26.098 50.322 26.181 ;
        RECT 44.802 14.69 110 15.5 ;
        RECT 50.276 9.216 50.322 26.181 ;
        RECT 33.348 26.144 50.276 26.227 ;
        RECT 44.848 14.644 110 15.5 ;
        RECT 50.23 9.262 50.276 26.227 ;
        RECT 33.302 26.19 50.23 26.273 ;
        RECT 44.894 14.598 110 15.5 ;
        RECT 50.184 9.308 50.23 26.273 ;
        RECT 33.256 26.236 50.184 26.319 ;
        RECT 44.94 14.552 110 15.5 ;
        RECT 50.138 9.354 50.184 26.319 ;
        RECT 33.21 26.282 50.138 26.365 ;
        RECT 44.986 14.506 110 15.5 ;
        RECT 50.092 9.4 50.138 26.365 ;
        RECT 33.164 26.328 50.092 26.411 ;
        RECT 45.032 14.46 110 15.5 ;
        RECT 50.046 9.446 50.092 26.411 ;
        RECT 33.118 26.374 50.046 26.457 ;
        RECT 45.078 14.414 110 15.5 ;
        RECT 50 9.492 50.046 26.457 ;
        RECT 33.072 26.42 50 26.503 ;
        RECT 45.124 14.368 110 15.5 ;
        RECT 49.954 9.538 50 26.503 ;
        RECT 33.026 26.466 49.954 26.549 ;
        RECT 45.17 14.322 110 15.5 ;
        RECT 49.908 9.584 49.954 26.549 ;
        RECT 32.98 26.512 49.908 26.595 ;
        RECT 45.216 14.276 110 15.5 ;
        RECT 49.862 9.63 49.908 26.595 ;
        RECT 32.934 26.558 49.862 26.641 ;
        RECT 45.262 14.23 110 15.5 ;
        RECT 49.816 9.676 49.862 26.641 ;
        RECT 32.888 26.604 49.816 26.687 ;
        RECT 45.308 14.184 110 15.5 ;
        RECT 49.77 9.722 49.816 26.687 ;
        RECT 32.842 26.65 49.77 26.733 ;
        RECT 45.354 14.138 110 15.5 ;
        RECT 49.724 9.768 49.77 26.733 ;
        RECT 32.796 26.696 49.724 26.779 ;
        RECT 45.4 14.092 110 15.5 ;
        RECT 49.678 9.814 49.724 26.779 ;
        RECT 32.75 26.742 49.678 26.825 ;
        RECT 45.446 14.046 110 15.5 ;
        RECT 49.632 9.86 49.678 26.825 ;
        RECT 32.704 26.788 49.632 26.871 ;
        RECT 45.492 14 110 15.5 ;
        RECT 49.586 9.906 49.632 26.871 ;
        RECT 32.658 26.834 49.586 26.917 ;
        RECT 45.538 13.954 110 15.5 ;
        RECT 49.54 9.952 49.586 26.917 ;
        RECT 32.612 26.88 49.54 26.963 ;
        RECT 45.584 13.908 110 15.5 ;
        RECT 49.494 9.998 49.54 26.963 ;
        RECT 32.566 26.926 49.494 27.009 ;
        RECT 45.63 13.862 110 15.5 ;
        RECT 49.448 10.044 49.494 27.009 ;
        RECT 32.52 26.972 49.448 27.055 ;
        RECT 45.676 13.816 110 15.5 ;
        RECT 49.402 10.09 49.448 27.055 ;
        RECT 32.474 27.018 49.402 27.101 ;
        RECT 45.722 13.77 110 15.5 ;
        RECT 49.356 10.136 49.402 27.101 ;
        RECT 32.428 27.064 49.356 27.147 ;
        RECT 45.768 13.724 110 15.5 ;
        RECT 49.31 10.182 49.356 27.147 ;
        RECT 32.382 27.11 49.31 27.193 ;
        RECT 45.814 13.678 110 15.5 ;
        RECT 49.264 10.228 49.31 27.193 ;
        RECT 32.336 27.156 49.264 27.239 ;
        RECT 45.86 13.632 110 15.5 ;
        RECT 49.218 10.274 49.264 27.239 ;
        RECT 32.29 27.202 49.218 27.285 ;
        RECT 45.906 13.586 110 15.5 ;
        RECT 49.172 10.32 49.218 27.285 ;
        RECT 32.244 27.248 49.172 27.331 ;
        RECT 45.952 13.54 110 15.5 ;
        RECT 49.126 10.366 49.172 27.331 ;
        RECT 32.198 27.294 49.126 27.377 ;
        RECT 45.998 13.494 110 15.5 ;
        RECT 49.08 10.412 49.126 27.377 ;
        RECT 32.152 27.34 49.08 27.423 ;
        RECT 46.044 13.448 110 15.5 ;
        RECT 49.034 10.458 49.08 27.423 ;
        RECT 32.106 27.386 49.034 27.469 ;
        RECT 46.09 13.402 110 15.5 ;
        RECT 48.988 10.504 49.034 27.469 ;
        RECT 32.06 27.432 48.988 27.515 ;
        RECT 46.136 13.356 110 15.5 ;
        RECT 48.942 10.55 48.988 27.515 ;
        RECT 32.014 27.478 48.942 27.561 ;
        RECT 46.182 13.31 110 15.5 ;
        RECT 48.896 10.596 48.942 27.561 ;
        RECT 31.968 27.524 48.896 27.607 ;
        RECT 46.228 13.264 110 15.5 ;
        RECT 48.85 10.642 48.896 27.607 ;
        RECT 31.922 27.57 48.85 27.653 ;
        RECT 46.274 13.218 110 15.5 ;
        RECT 48.804 10.688 48.85 27.653 ;
        RECT 31.876 27.616 48.804 27.699 ;
        RECT 46.32 13.172 110 15.5 ;
        RECT 48.758 10.734 48.804 27.699 ;
        RECT 31.83 27.662 48.758 27.745 ;
        RECT 46.366 13.126 110 15.5 ;
        RECT 48.712 10.78 48.758 27.745 ;
        RECT 31.784 27.708 48.712 27.791 ;
        RECT 46.412 13.08 110 15.5 ;
        RECT 48.666 10.826 48.712 27.791 ;
        RECT 31.738 27.754 48.666 27.837 ;
        RECT 46.458 13.034 110 15.5 ;
        RECT 48.62 10.872 48.666 27.837 ;
        RECT 31.692 27.8 48.62 27.883 ;
        RECT 46.504 12.988 110 15.5 ;
        RECT 48.574 10.918 48.62 27.883 ;
        RECT 31.646 27.846 48.574 27.929 ;
        RECT 46.55 12.942 110 15.5 ;
        RECT 48.528 10.964 48.574 27.929 ;
        RECT 31.6 27.892 48.528 27.975 ;
        RECT 46.596 12.896 110 15.5 ;
        RECT 48.482 11.01 48.528 27.975 ;
        RECT 31.554 27.938 48.482 28.021 ;
        RECT 46.642 12.85 110 15.5 ;
        RECT 48.436 11.056 48.482 28.021 ;
        RECT 31.508 27.984 48.436 28.067 ;
        RECT 46.688 12.804 110 15.5 ;
        RECT 48.39 11.102 48.436 28.067 ;
        RECT 31.462 28.03 48.39 28.113 ;
        RECT 46.734 12.758 110 15.5 ;
        RECT 48.344 11.148 48.39 28.113 ;
        RECT 31.416 28.076 48.344 28.159 ;
        RECT 46.78 12.712 110 15.5 ;
        RECT 48.298 11.194 48.344 28.159 ;
        RECT 31.37 28.122 48.298 28.205 ;
        RECT 46.826 12.666 110 15.5 ;
        RECT 48.252 11.24 48.298 28.205 ;
        RECT 31.324 28.168 48.252 28.251 ;
        RECT 46.872 12.62 110 15.5 ;
        RECT 48.206 11.286 48.252 28.251 ;
        RECT 31.278 28.214 48.206 28.297 ;
        RECT 46.918 12.574 110 15.5 ;
        RECT 48.16 11.332 48.206 28.297 ;
        RECT 31.232 28.26 48.16 28.343 ;
        RECT 46.964 12.528 110 15.5 ;
        RECT 48.114 11.378 48.16 28.343 ;
        RECT 31.186 28.306 48.114 28.389 ;
        RECT 47.01 12.482 110 15.5 ;
        RECT 48.068 11.424 48.114 28.389 ;
        RECT 31.14 28.352 48.068 28.435 ;
        RECT 47.056 12.436 110 15.5 ;
        RECT 48.022 11.47 48.068 28.435 ;
        RECT 31.094 28.398 48.022 28.481 ;
        RECT 47.102 12.39 110 15.5 ;
        RECT 47.976 11.516 48.022 28.481 ;
        RECT 31.048 28.444 47.976 28.527 ;
        RECT 47.148 12.344 110 15.5 ;
        RECT 47.93 11.562 47.976 28.527 ;
        RECT 31.002 28.49 47.93 28.573 ;
        RECT 47.194 12.298 110 15.5 ;
        RECT 47.884 11.608 47.93 28.573 ;
        RECT 30.956 28.536 47.884 28.619 ;
        RECT 47.24 12.252 110 15.5 ;
        RECT 47.838 11.654 47.884 28.619 ;
        RECT 30.91 28.582 47.838 28.665 ;
        RECT 47.286 12.206 110 15.5 ;
        RECT 47.792 11.7 47.838 28.665 ;
        RECT 30.864 28.628 47.792 28.711 ;
        RECT 47.332 12.16 110 15.5 ;
        RECT 47.746 11.746 47.792 28.711 ;
        RECT 30.818 28.674 47.746 28.757 ;
        RECT 47.378 12.114 110 15.5 ;
        RECT 47.7 11.792 47.746 28.757 ;
        RECT 30.772 28.72 47.7 28.803 ;
        RECT 47.424 12.068 110 15.5 ;
        RECT 47.654 11.838 47.7 28.803 ;
        RECT 30.726 28.766 47.654 28.849 ;
        RECT 47.47 12.022 110 15.5 ;
        RECT 47.608 11.884 47.654 28.849 ;
        RECT 30.68 28.812 47.608 28.895 ;
        RECT 47.516 11.976 110 15.5 ;
        RECT 47.562 11.93 47.608 28.895 ;
        RECT 30.634 28.858 47.562 28.941 ;
        RECT 30.588 28.904 47.516 28.987 ;
        RECT 30.542 28.95 47.47 29.033 ;
        RECT 30.496 28.996 47.424 29.079 ;
        RECT 30.45 29.042 47.378 29.125 ;
        RECT 30.404 29.088 47.332 29.171 ;
        RECT 30.358 29.134 47.286 29.217 ;
        RECT 30.312 29.18 47.24 29.263 ;
        RECT 30.266 29.226 47.194 29.309 ;
        RECT 30.22 29.272 47.148 29.355 ;
        RECT 30.174 29.318 47.102 29.401 ;
        RECT 30.128 29.364 47.056 29.447 ;
        RECT 30.082 29.41 47.01 29.493 ;
        RECT 30.036 29.456 46.964 29.539 ;
        RECT 29.99 29.502 46.918 29.585 ;
        RECT 29.944 29.548 46.872 29.631 ;
        RECT 29.898 29.594 46.826 29.677 ;
        RECT 29.852 29.64 46.78 29.723 ;
        RECT 29.806 29.686 46.734 29.769 ;
        RECT 29.76 29.732 46.688 29.815 ;
        RECT 29.714 29.778 46.642 29.861 ;
        RECT 29.668 29.824 46.596 29.907 ;
        RECT 29.622 29.87 46.55 29.953 ;
        RECT 29.576 29.916 46.504 29.999 ;
        RECT 29.53 29.962 46.458 30.045 ;
        RECT 29.484 30.008 46.412 30.091 ;
        RECT 29.438 30.054 46.366 30.137 ;
        RECT 29.392 30.1 46.32 30.183 ;
        RECT 29.346 30.146 46.274 30.229 ;
        RECT 29.3 30.192 46.228 30.275 ;
        RECT 29.254 30.238 46.182 30.321 ;
        RECT 29.208 30.284 46.136 30.367 ;
        RECT 29.162 30.33 46.09 30.413 ;
        RECT 29.116 30.376 46.044 30.459 ;
        RECT 29.07 30.422 45.998 30.505 ;
        RECT 29.024 30.468 45.952 30.551 ;
        RECT 28.978 30.514 45.906 30.597 ;
        RECT 28.932 30.56 45.86 30.643 ;
        RECT 28.886 30.606 45.814 30.689 ;
        RECT 28.84 30.652 45.768 30.735 ;
        RECT 28.794 30.698 45.722 30.781 ;
        RECT 28.748 30.744 45.676 30.827 ;
        RECT 28.702 30.79 45.63 30.873 ;
        RECT 28.656 30.836 45.584 30.919 ;
        RECT 28.61 30.882 45.538 30.965 ;
        RECT 28.564 30.928 45.492 31.011 ;
        RECT 28.518 30.974 45.446 31.057 ;
        RECT 28.472 31.02 45.4 31.103 ;
        RECT 28.426 31.066 45.354 31.149 ;
        RECT 28.38 31.112 45.308 31.195 ;
        RECT 28.334 31.158 45.262 31.241 ;
        RECT 28.288 31.204 45.216 31.287 ;
        RECT 28.242 31.25 45.17 31.333 ;
        RECT 28.196 31.296 45.124 31.379 ;
        RECT 28.15 31.342 45.078 31.425 ;
        RECT 28.104 31.388 45.032 31.471 ;
        RECT 28.058 31.434 44.986 31.517 ;
        RECT 28.012 31.48 44.94 31.563 ;
        RECT 27.966 31.526 44.894 31.609 ;
        RECT 27.92 31.572 44.848 31.655 ;
        RECT 27.874 31.618 44.802 31.701 ;
        RECT 27.828 31.664 44.756 31.747 ;
        RECT 27.782 31.71 44.71 31.793 ;
        RECT 27.736 31.756 44.664 31.839 ;
        RECT 27.69 31.802 44.618 31.885 ;
        RECT 27.644 31.848 44.572 31.931 ;
        RECT 27.598 31.894 44.526 31.977 ;
        RECT 27.552 31.94 44.48 32.023 ;
        RECT 27.506 31.986 44.434 32.069 ;
        RECT 27.46 32.032 44.388 32.115 ;
        RECT 27.414 32.078 44.342 32.161 ;
        RECT 27.368 32.124 44.296 32.207 ;
        RECT 27.322 32.17 44.25 32.253 ;
        RECT 27.276 32.216 44.204 32.299 ;
        RECT 27.23 32.262 44.158 32.345 ;
        RECT 27.184 32.308 44.112 32.391 ;
        RECT 27.138 32.354 44.066 32.437 ;
        RECT 27.092 32.4 44.02 32.483 ;
        RECT 27.046 32.446 43.974 32.529 ;
        RECT 27 32.492 43.928 32.575 ;
        RECT 26.954 32.538 43.882 32.621 ;
        RECT 26.908 32.584 43.836 32.667 ;
        RECT 26.862 32.63 43.79 32.713 ;
        RECT 26.816 32.676 43.744 32.759 ;
        RECT 26.77 32.722 43.698 32.805 ;
        RECT 26.724 32.768 43.652 32.851 ;
        RECT 26.678 32.814 43.606 32.897 ;
        RECT 26.632 32.86 43.56 32.943 ;
        RECT 26.586 32.906 43.514 32.989 ;
        RECT 26.54 32.952 43.468 33.035 ;
        RECT 26.494 32.998 43.422 33.081 ;
        RECT 26.448 33.044 43.376 33.127 ;
        RECT 26.402 33.09 43.33 33.173 ;
        RECT 26.356 33.136 43.284 33.219 ;
        RECT 26.31 33.182 43.238 33.265 ;
        RECT 26.264 33.228 43.192 33.311 ;
        RECT 26.218 33.274 43.146 33.357 ;
        RECT 26.172 33.32 43.1 33.403 ;
        RECT 26.126 33.366 43.054 33.449 ;
        RECT 26.08 33.412 43.008 33.495 ;
        RECT 26.034 33.458 42.962 33.541 ;
        RECT 25.988 33.504 42.916 33.587 ;
        RECT 25.942 33.55 42.87 33.633 ;
        RECT 25.896 33.596 42.824 33.679 ;
        RECT 25.85 33.642 42.778 33.725 ;
        RECT 25.804 33.688 42.732 33.771 ;
        RECT 25.758 33.734 42.686 33.817 ;
        RECT 25.712 33.78 42.64 33.863 ;
        RECT 25.666 33.826 42.594 33.909 ;
        RECT 25.62 33.872 42.548 33.955 ;
        RECT 25.574 33.918 42.502 34.001 ;
        RECT 25.528 33.964 42.456 34.047 ;
        RECT 25.482 34.01 42.41 34.093 ;
        RECT 25.436 34.056 42.364 34.139 ;
        RECT 25.39 34.102 42.318 34.185 ;
        RECT 25.344 34.148 42.272 34.231 ;
        RECT 25.298 34.194 42.226 34.277 ;
        RECT 25.252 34.24 42.18 34.323 ;
        RECT 25.206 34.286 42.134 34.369 ;
        RECT 25.16 34.332 42.088 34.415 ;
        RECT 25.114 34.378 42.042 34.461 ;
        RECT 25.068 34.424 41.996 34.507 ;
        RECT 25.022 34.47 41.95 34.553 ;
        RECT 24.976 34.516 41.904 34.599 ;
        RECT 24.93 34.562 41.858 34.645 ;
        RECT 24.884 34.608 41.812 34.691 ;
        RECT 24.838 34.654 41.766 34.737 ;
        RECT 24.792 34.7 41.72 34.783 ;
        RECT 24.746 34.746 41.674 34.829 ;
        RECT 24.7 34.792 41.628 34.875 ;
        RECT 24.654 34.838 41.582 34.921 ;
        RECT 24.608 34.884 41.536 34.967 ;
        RECT 24.562 34.93 41.49 35.013 ;
        RECT 24.516 34.976 41.444 35.059 ;
        RECT 24.47 35.022 41.398 35.105 ;
        RECT 24.424 35.068 41.352 35.151 ;
        RECT 24.378 35.114 41.306 35.197 ;
        RECT 24.332 35.16 41.26 35.243 ;
        RECT 24.286 35.206 41.214 35.289 ;
        RECT 24.24 35.252 41.168 35.335 ;
        RECT 24.194 35.298 41.122 35.381 ;
        RECT 24.148 35.344 41.076 35.427 ;
        RECT 24.102 35.39 41.03 35.473 ;
        RECT 24.056 35.436 40.984 35.519 ;
        RECT 24.01 35.482 40.938 35.565 ;
        RECT 23.964 35.528 40.892 35.611 ;
        RECT 23.918 35.574 40.846 35.657 ;
        RECT 23.872 35.62 40.8 35.703 ;
        RECT 23.826 35.666 40.754 35.749 ;
        RECT 23.78 35.712 40.708 35.795 ;
        RECT 23.734 35.758 40.662 35.841 ;
        RECT 23.688 35.804 40.616 35.887 ;
        RECT 23.642 35.85 40.57 35.933 ;
        RECT 23.596 35.896 40.524 35.979 ;
        RECT 23.55 35.942 40.478 36.025 ;
        RECT 23.504 35.988 40.432 36.071 ;
        RECT 23.458 36.034 40.386 36.117 ;
        RECT 23.412 36.08 40.34 36.163 ;
        RECT 23.366 36.126 40.294 36.209 ;
        RECT 23.32 36.172 40.248 36.255 ;
        RECT 23.274 36.218 40.202 36.301 ;
        RECT 23.228 36.264 40.156 36.347 ;
        RECT 23.182 36.31 40.11 36.393 ;
        RECT 23.136 36.356 40.064 36.439 ;
        RECT 23.09 36.402 40.018 36.485 ;
        RECT 23.044 36.448 39.972 36.531 ;
        RECT 22.998 36.494 39.926 36.577 ;
        RECT 22.952 36.54 39.88 36.623 ;
        RECT 22.906 36.586 39.834 36.669 ;
        RECT 22.86 36.632 39.788 36.715 ;
        RECT 22.814 36.678 39.742 36.761 ;
        RECT 22.768 36.724 39.696 36.807 ;
        RECT 22.722 36.77 39.65 36.853 ;
        RECT 22.676 36.816 39.604 36.899 ;
        RECT 22.63 36.862 39.558 36.945 ;
        RECT 22.584 36.908 39.512 36.991 ;
        RECT 22.538 36.954 39.466 37.037 ;
        RECT 22.492 37 39.42 37.083 ;
        RECT 22.446 37.046 39.374 37.129 ;
        RECT 22.4 37.092 39.328 37.175 ;
        RECT 22.354 37.138 39.282 37.221 ;
        RECT 22.308 37.184 39.236 37.267 ;
        RECT 22.262 37.23 39.19 37.313 ;
        RECT 22.216 37.276 39.144 37.359 ;
        RECT 22.17 37.322 39.098 37.405 ;
        RECT 22.124 37.368 39.052 37.451 ;
        RECT 22.078 37.414 39.006 37.497 ;
        RECT 22.032 37.46 38.96 37.543 ;
        RECT 21.986 37.506 38.914 37.589 ;
        RECT 21.94 37.552 38.868 37.635 ;
        RECT 21.894 37.598 38.822 37.681 ;
        RECT 21.848 37.644 38.776 37.727 ;
        RECT 21.802 37.69 38.73 37.773 ;
        RECT 21.756 37.736 38.684 37.819 ;
        RECT 21.71 37.782 38.638 37.865 ;
        RECT 21.664 37.828 38.592 37.911 ;
        RECT 21.618 37.874 38.546 37.957 ;
        RECT 21.572 37.92 38.5 38.003 ;
        RECT 21.526 37.966 38.454 38.049 ;
        RECT 21.48 38.012 38.408 38.095 ;
        RECT 21.434 38.058 38.362 38.141 ;
        RECT 21.388 38.104 38.316 38.187 ;
        RECT 21.342 38.15 38.27 38.233 ;
        RECT 21.296 38.196 38.224 38.279 ;
        RECT 21.25 38.242 38.178 38.325 ;
        RECT 21.204 38.288 38.132 38.371 ;
        RECT 21.158 38.334 38.086 38.417 ;
        RECT 21.112 38.38 38.04 38.463 ;
        RECT 21.066 38.426 37.994 38.509 ;
        RECT 21.02 38.472 37.948 38.555 ;
        RECT 20.974 38.518 37.902 38.601 ;
        RECT 20.928 38.564 37.856 38.647 ;
        RECT 20.882 38.61 37.81 38.693 ;
        RECT 20.836 38.656 37.764 38.739 ;
        RECT 20.79 38.702 37.718 38.785 ;
        RECT 20.744 38.748 37.672 38.831 ;
        RECT 20.698 38.794 37.626 38.877 ;
        RECT 20.652 38.84 37.58 38.923 ;
        RECT 20.606 38.886 37.534 38.969 ;
        RECT 20.56 38.932 37.488 39.015 ;
        RECT 20.514 38.978 37.442 39.061 ;
        RECT 20.468 39.024 37.396 39.107 ;
        RECT 20.422 39.07 37.35 39.153 ;
        RECT 20.376 39.116 37.304 39.199 ;
        RECT 20.33 39.162 37.258 39.245 ;
        RECT 20.284 39.208 37.212 39.291 ;
        RECT 20.238 39.254 37.166 39.337 ;
        RECT 20.192 39.3 37.12 39.383 ;
        RECT 20.146 39.346 37.074 39.429 ;
        RECT 20.1 39.392 37.028 39.475 ;
        RECT 20.054 39.438 36.982 39.521 ;
        RECT 20.008 39.484 36.936 39.567 ;
        RECT 19.962 39.53 36.89 39.613 ;
        RECT 19.916 39.576 36.844 39.659 ;
        RECT 19.87 39.622 36.798 39.705 ;
        RECT 19.824 39.668 36.752 39.751 ;
        RECT 19.778 39.714 36.706 39.797 ;
        RECT 19.732 39.76 36.66 39.843 ;
        RECT 19.686 39.806 36.614 39.889 ;
        RECT 19.64 39.852 36.568 39.935 ;
        RECT 19.594 39.898 36.522 39.981 ;
        RECT 19.548 39.944 36.476 40.027 ;
        RECT 19.502 39.99 36.43 40.073 ;
        RECT 19.456 40.036 36.384 40.119 ;
        RECT 19.41 40.082 36.338 40.165 ;
        RECT 19.364 40.128 36.292 40.211 ;
        RECT 19.318 40.174 36.246 40.257 ;
        RECT 19.272 40.22 36.2 40.303 ;
        RECT 19.226 40.266 36.154 40.349 ;
        RECT 19.18 40.312 36.108 40.395 ;
        RECT 19.134 40.358 36.062 40.441 ;
        RECT 19.088 40.404 36.016 40.487 ;
        RECT 19.042 40.45 35.97 40.533 ;
        RECT 18.996 40.496 35.924 40.579 ;
        RECT 18.95 40.542 35.878 40.625 ;
        RECT 18.904 40.588 35.832 40.671 ;
        RECT 18.858 40.634 35.786 40.717 ;
        RECT 18.812 40.68 35.74 40.763 ;
        RECT 18.766 40.726 35.694 40.809 ;
        RECT 18.72 40.772 35.648 40.855 ;
        RECT 18.674 40.818 35.602 40.901 ;
        RECT 18.628 40.864 35.556 40.947 ;
        RECT 18.582 40.91 35.51 40.993 ;
        RECT 18.536 40.956 35.464 41.039 ;
        RECT 18.49 41.002 35.418 41.085 ;
        RECT 18.444 41.048 35.372 41.131 ;
        RECT 18.398 41.094 35.326 41.177 ;
        RECT 18.352 41.14 35.28 41.223 ;
        RECT 18.306 41.186 35.234 41.269 ;
        RECT 18.26 41.232 35.188 41.315 ;
        RECT 18.214 41.278 35.142 41.361 ;
        RECT 18.168 41.324 35.096 41.407 ;
        RECT 18.122 41.37 35.05 41.453 ;
        RECT 18.076 41.416 35.004 41.499 ;
        RECT 18.03 41.462 34.958 41.545 ;
        RECT 17.984 41.508 34.912 41.591 ;
        RECT 17.938 41.554 34.866 41.637 ;
        RECT 17.892 41.6 34.82 41.683 ;
        RECT 17.846 41.646 34.774 41.729 ;
        RECT 17.8 41.692 34.728 41.775 ;
        RECT 17.754 41.738 34.682 41.821 ;
        RECT 17.708 41.784 34.636 41.867 ;
        RECT 17.662 41.83 34.59 41.913 ;
        RECT 17.616 41.876 34.544 41.959 ;
        RECT 17.57 41.922 34.498 42.005 ;
        RECT 17.524 41.968 34.452 42.051 ;
        RECT 17.478 42.014 34.406 42.097 ;
        RECT 17.432 42.06 34.36 42.143 ;
        RECT 17.386 42.106 34.314 42.189 ;
        RECT 17.34 42.152 34.268 42.235 ;
        RECT 17.294 42.198 34.222 42.281 ;
        RECT 17.248 42.244 34.176 42.327 ;
        RECT 17.202 42.29 34.13 42.373 ;
        RECT 17.156 42.336 34.084 42.419 ;
        RECT 17.11 42.382 34.038 42.465 ;
        RECT 17.064 42.428 33.992 42.511 ;
        RECT 17.018 42.474 33.946 42.557 ;
        RECT 16.972 42.52 33.9 42.603 ;
        RECT 16.926 42.566 33.854 42.649 ;
        RECT 16.88 42.612 33.808 42.695 ;
        RECT 16.834 42.658 33.762 42.741 ;
        RECT 16.788 42.704 33.716 42.787 ;
        RECT 16.742 42.75 33.67 42.833 ;
        RECT 16.696 42.796 33.624 42.879 ;
        RECT 16.65 42.842 33.578 42.925 ;
        RECT 16.604 42.888 33.532 42.971 ;
        RECT 16.558 42.934 33.486 43.017 ;
        RECT 16.512 42.98 33.44 43.063 ;
        RECT 16.466 43.026 33.394 43.109 ;
        RECT 16.42 43.072 33.348 43.155 ;
        RECT 16.374 43.118 33.302 43.201 ;
        RECT 16.328 43.164 33.256 43.247 ;
        RECT 16.282 43.21 33.21 43.293 ;
        RECT 16.236 43.256 33.164 43.339 ;
        RECT 16.19 43.302 33.118 43.385 ;
        RECT 16.144 43.348 33.072 43.431 ;
        RECT 16.098 43.394 33.026 43.477 ;
        RECT 16.052 43.44 32.98 43.523 ;
        RECT 16.006 43.486 32.934 43.569 ;
        RECT 15.96 43.532 32.888 43.615 ;
        RECT 15.914 43.578 32.842 43.661 ;
        RECT 15.868 43.624 32.796 43.707 ;
        RECT 15.822 43.67 32.75 43.753 ;
        RECT 15.776 43.716 32.704 43.799 ;
        RECT 15.73 43.762 32.658 43.845 ;
        RECT 15.684 43.808 32.612 43.891 ;
        RECT 15.638 43.854 32.566 43.937 ;
        RECT 15.592 43.9 32.52 43.983 ;
        RECT 15.546 43.946 32.474 44.029 ;
        RECT 15.5 43.992 32.428 44.075 ;
        RECT 15.46 44.035 32.382 44.121 ;
        RECT 15.414 44.078 32.336 44.167 ;
        RECT 15.368 44.124 32.29 44.213 ;
        RECT 15.322 44.17 32.244 44.259 ;
        RECT 15.276 44.216 32.198 44.305 ;
        RECT 15.23 44.262 32.152 44.351 ;
        RECT 15.184 44.308 32.106 44.397 ;
        RECT 15.138 44.354 32.06 44.443 ;
        RECT 15.092 44.4 32.014 44.489 ;
        RECT 15.046 44.446 31.968 44.535 ;
        RECT 15 44.492 31.922 44.581 ;
        RECT 14.954 44.538 31.876 44.627 ;
        RECT 14.908 44.584 31.83 44.673 ;
        RECT 14.862 44.63 31.784 44.719 ;
        RECT 14.816 44.676 31.738 44.765 ;
        RECT 14.77 44.722 31.692 44.811 ;
        RECT 14.724 44.768 31.646 44.857 ;
        RECT 14.678 44.814 31.6 44.903 ;
        RECT 14.632 44.86 31.554 44.949 ;
        RECT 14.586 44.906 31.508 44.995 ;
        RECT 14.54 44.952 31.462 45.041 ;
        RECT 14.494 44.998 31.416 45.087 ;
        RECT 14.448 45.044 31.37 45.133 ;
        RECT 14.402 45.09 31.324 45.179 ;
        RECT 14.356 45.136 31.278 45.225 ;
        RECT 14.31 45.182 31.232 45.271 ;
        RECT 14.264 45.228 31.186 45.317 ;
        RECT 14.218 45.274 31.14 45.363 ;
        RECT 14.172 45.32 31.094 45.409 ;
        RECT 14.126 45.366 31.048 45.455 ;
        RECT 14.08 45.412 31.002 45.501 ;
        RECT 14.034 45.458 30.956 45.547 ;
        RECT 13.988 45.504 30.91 45.593 ;
        RECT 13.942 45.55 30.864 45.639 ;
        RECT 13.896 45.596 30.818 45.685 ;
        RECT 13.85 45.642 30.772 45.731 ;
        RECT 13.804 45.688 30.726 45.777 ;
        RECT 13.758 45.734 30.68 45.823 ;
        RECT 13.712 45.78 30.634 45.869 ;
        RECT 13.666 45.826 30.588 45.915 ;
        RECT 13.62 45.872 30.542 45.961 ;
        RECT 13.574 45.918 30.496 46.007 ;
        RECT 13.528 45.964 30.45 46.053 ;
        RECT 13.482 46.01 30.404 46.099 ;
        RECT 13.436 46.056 30.358 46.145 ;
        RECT 13.39 46.102 30.312 46.191 ;
        RECT 13.344 46.148 30.266 46.237 ;
        RECT 13.298 46.194 30.22 46.283 ;
        RECT 13.252 46.24 30.174 46.329 ;
        RECT 13.206 46.286 30.128 46.375 ;
        RECT 13.16 46.332 30.082 46.421 ;
        RECT 13.114 46.378 30.036 46.467 ;
        RECT 13.068 46.424 29.99 46.513 ;
        RECT 13.022 46.47 29.944 46.559 ;
        RECT 12.976 46.516 29.898 46.605 ;
        RECT 12.93 46.562 29.852 46.651 ;
        RECT 12.884 46.608 29.806 46.697 ;
        RECT 12.838 46.654 29.76 46.743 ;
        RECT 12.792 46.7 29.714 46.789 ;
        RECT 12.746 46.746 29.668 46.835 ;
        RECT 12.7 46.792 29.622 46.881 ;
        RECT 12.654 46.838 29.576 46.927 ;
        RECT 12.608 46.884 29.53 46.973 ;
        RECT 12.562 46.93 29.484 47.019 ;
        RECT 12.516 46.976 29.438 47.065 ;
        RECT 12.47 47.022 29.392 47.111 ;
        RECT 12.424 47.068 29.346 47.157 ;
        RECT 12.378 47.114 29.3 47.203 ;
        RECT 12.332 47.16 29.254 47.249 ;
        RECT 12.286 47.206 29.208 47.295 ;
        RECT 12.24 47.252 29.162 47.341 ;
        RECT 12.194 47.298 29.116 47.387 ;
        RECT 12.148 47.344 29.07 47.433 ;
        RECT 12.102 47.39 29.024 47.479 ;
        RECT 12.056 47.436 28.978 47.525 ;
        RECT 12.01 47.482 28.932 47.571 ;
        RECT 11.964 47.528 28.886 47.617 ;
        RECT 11.918 47.574 28.84 47.663 ;
        RECT 11.872 47.62 28.794 47.709 ;
        RECT 11.826 47.666 28.748 47.755 ;
        RECT 11.78 47.712 28.702 47.801 ;
        RECT 11.734 47.758 28.656 47.847 ;
        RECT 11.688 47.804 28.61 47.893 ;
        RECT 11.642 47.85 28.564 47.939 ;
        RECT 11.596 47.896 28.518 47.985 ;
        RECT 11.55 47.942 28.472 48.031 ;
        RECT 11.504 47.988 28.426 48.077 ;
        RECT 11.458 48.034 28.38 48.123 ;
        RECT 11.412 48.08 28.334 48.169 ;
        RECT 11.366 48.126 28.288 48.215 ;
        RECT 11.32 48.172 28.242 48.261 ;
        RECT 11.274 48.218 28.196 48.307 ;
        RECT 11.228 48.264 28.15 48.353 ;
        RECT 11.182 48.31 28.104 48.399 ;
        RECT 11.136 48.356 28.058 48.445 ;
        RECT 11.09 48.402 28.012 48.491 ;
        RECT 11.044 48.448 27.966 48.537 ;
        RECT 10.998 48.494 27.92 48.583 ;
        RECT 10.952 48.54 27.874 48.629 ;
        RECT 10.906 48.586 27.828 48.675 ;
        RECT 10.86 48.632 27.782 48.721 ;
        RECT 10.814 48.678 27.736 48.767 ;
        RECT 10.768 48.724 27.69 48.813 ;
        RECT 10.722 48.77 27.644 48.859 ;
        RECT 10.676 48.816 27.598 48.905 ;
        RECT 10.63 48.862 27.552 48.951 ;
        RECT 10.584 48.908 27.506 48.997 ;
        RECT 10.538 48.954 27.46 49.043 ;
        RECT 10.492 49 27.414 49.089 ;
        RECT 10.446 49.046 27.368 49.135 ;
        RECT 10.4 49.092 27.322 49.181 ;
        RECT 10.354 49.138 27.276 49.227 ;
        RECT 10.308 49.184 27.23 49.273 ;
        RECT 10.262 49.23 27.184 49.319 ;
        RECT 10.216 49.276 27.138 49.365 ;
        RECT 10.17 49.322 27.092 49.411 ;
        RECT 10.124 49.368 27.046 49.457 ;
        RECT 10.078 49.414 27 49.503 ;
      LAYER MET4 ;
        RECT 28.362 51.38 45.33 51.428 ;
        RECT 28.316 51.426 45.284 51.474 ;
        RECT 28.27 51.472 45.238 51.52 ;
        RECT 28.224 51.518 45.192 51.566 ;
        RECT 28.178 51.564 45.146 51.612 ;
        RECT 28.132 51.61 45.1 51.658 ;
        RECT 28.086 51.656 45.054 51.704 ;
        RECT 28.04 51.702 45.008 51.75 ;
        RECT 27.994 51.748 44.962 51.796 ;
        RECT 27.948 51.794 44.916 51.842 ;
        RECT 27.902 51.84 44.87 51.888 ;
        RECT 27.856 51.886 44.824 51.934 ;
        RECT 27.81 51.932 44.778 51.98 ;
        RECT 27.764 51.978 44.732 52.026 ;
        RECT 27.718 52.024 44.686 52.072 ;
        RECT 27.672 52.07 44.64 52.118 ;
        RECT 27.626 52.116 44.594 52.164 ;
        RECT 27.58 52.162 44.548 52.21 ;
        RECT 27.534 52.208 44.502 52.256 ;
        RECT 27.488 52.254 44.456 52.302 ;
        RECT 27.442 52.3 44.41 52.348 ;
        RECT 27.396 52.346 44.364 52.394 ;
        RECT 27.35 52.392 44.318 52.44 ;
        RECT 27.304 52.438 44.272 52.486 ;
        RECT 27.258 52.484 44.226 52.532 ;
        RECT 27.212 52.53 44.18 52.578 ;
        RECT 27.166 52.576 44.134 52.624 ;
        RECT 27.12 52.622 44.088 52.67 ;
        RECT 27.074 52.668 44.042 52.716 ;
        RECT 27.028 52.714 43.996 52.762 ;
        RECT 26.982 52.76 43.95 52.808 ;
        RECT 26.936 52.806 43.904 52.854 ;
        RECT 26.89 52.852 43.858 52.9 ;
        RECT 26.844 52.898 43.812 52.946 ;
        RECT 26.798 52.944 43.766 52.992 ;
        RECT 26.752 52.99 43.72 53.038 ;
        RECT 26.706 53.036 43.674 53.084 ;
        RECT 26.66 53.082 43.628 53.13 ;
        RECT 26.614 53.128 43.582 53.176 ;
        RECT 26.568 53.174 43.536 53.222 ;
        RECT 26.522 53.22 43.49 53.268 ;
        RECT 26.476 53.266 43.444 53.314 ;
        RECT 26.43 53.312 43.398 53.36 ;
        RECT 26.384 53.358 43.352 53.406 ;
        RECT 26.338 53.404 43.306 53.452 ;
        RECT 26.292 53.45 43.26 53.498 ;
        RECT 26.246 53.496 43.214 53.544 ;
        RECT 26.2 53.542 43.168 53.59 ;
        RECT 26.154 53.588 43.122 53.636 ;
        RECT 26.108 53.634 43.076 53.682 ;
        RECT 26.062 53.68 43.03 53.728 ;
        RECT 26.016 53.726 42.984 53.774 ;
        RECT 25.97 53.772 42.938 53.82 ;
        RECT 25.924 53.818 42.892 53.866 ;
        RECT 25.878 53.864 42.846 53.912 ;
        RECT 25.832 53.91 42.8 53.958 ;
        RECT 25.786 53.956 42.754 54.004 ;
        RECT 25.74 54.002 42.708 54.05 ;
        RECT 25.694 54.048 42.662 54.096 ;
        RECT 25.648 54.094 42.616 54.142 ;
        RECT 25.602 54.14 42.57 54.188 ;
        RECT 25.556 54.186 42.524 54.234 ;
        RECT 25.51 54.232 42.478 54.28 ;
        RECT 25.464 54.278 42.432 54.326 ;
        RECT 25.418 54.324 42.386 54.372 ;
        RECT 25.372 54.37 42.34 54.418 ;
        RECT 25.326 54.416 42.294 54.464 ;
        RECT 25.28 54.462 42.248 54.51 ;
        RECT 25.234 54.508 42.202 54.556 ;
        RECT 25.188 54.554 42.156 54.602 ;
        RECT 25.142 54.6 42.11 54.648 ;
        RECT 25.096 54.646 42.064 54.694 ;
        RECT 25.05 54.692 42.018 54.74 ;
        RECT 25.004 54.738 41.972 54.786 ;
        RECT 24.958 54.784 41.926 54.832 ;
        RECT 24.912 54.83 41.88 54.878 ;
        RECT 24.866 54.876 41.834 54.924 ;
        RECT 24.82 54.922 41.788 54.97 ;
        RECT 24.774 54.968 41.742 55.016 ;
        RECT 24.728 55.014 41.696 55.062 ;
        RECT 24.682 55.06 41.65 55.108 ;
        RECT 24.636 55.106 41.604 55.154 ;
        RECT 24.59 55.152 41.558 55.2 ;
        RECT 24.544 55.198 41.512 55.246 ;
        RECT 24.498 55.244 41.466 55.292 ;
        RECT 24.452 55.29 41.42 55.338 ;
        RECT 24.406 55.336 41.374 55.384 ;
        RECT 24.36 55.382 41.328 55.43 ;
        RECT 24.314 55.428 41.282 55.476 ;
        RECT 24.268 55.474 41.236 55.522 ;
        RECT 24.222 55.52 41.19 55.568 ;
        RECT 24.176 55.566 41.144 55.614 ;
        RECT 24.13 55.612 41.098 55.66 ;
        RECT 24.084 55.658 41.052 55.706 ;
        RECT 24.038 55.704 41.006 55.752 ;
        RECT 23.992 55.75 40.96 55.798 ;
        RECT 23.946 55.796 40.914 55.844 ;
        RECT 23.9 55.842 40.868 55.89 ;
        RECT 23.854 55.888 40.822 55.936 ;
        RECT 23.808 55.934 40.776 55.982 ;
        RECT 23.762 55.98 40.73 56.028 ;
        RECT 23.716 56.026 40.684 56.074 ;
        RECT 23.67 56.072 40.638 56.12 ;
        RECT 23.624 56.118 40.592 56.166 ;
        RECT 23.578 56.164 40.546 56.212 ;
        RECT 23.532 56.21 40.5 56.258 ;
        RECT 23.486 56.256 40.454 56.304 ;
        RECT 23.44 56.302 40.408 56.35 ;
        RECT 23.394 56.348 40.362 56.396 ;
        RECT 23.348 56.394 40.316 56.442 ;
        RECT 23.302 56.44 40.27 56.488 ;
        RECT 23.256 56.486 40.224 56.534 ;
        RECT 23.21 56.532 40.178 56.58 ;
        RECT 23.164 56.578 40.132 56.626 ;
        RECT 23.118 56.624 40.086 56.672 ;
        RECT 23.072 56.67 40.04 56.718 ;
        RECT 23.026 56.716 39.994 56.764 ;
        RECT 22.98 56.762 39.948 56.81 ;
        RECT 22.934 56.808 39.902 56.856 ;
        RECT 22.888 56.854 39.856 56.902 ;
        RECT 22.842 56.9 39.81 56.948 ;
        RECT 22.796 56.946 39.764 56.994 ;
        RECT 22.75 56.992 39.718 57.04 ;
        RECT 22.704 57.038 39.672 57.086 ;
        RECT 22.658 57.084 39.626 57.132 ;
        RECT 22.612 57.13 39.58 57.178 ;
        RECT 22.566 57.176 39.534 57.224 ;
        RECT 22.52 57.222 39.488 57.27 ;
        RECT 22.474 57.268 39.442 57.316 ;
        RECT 22.428 57.314 39.396 57.362 ;
        RECT 22.382 57.36 39.35 57.408 ;
        RECT 22.336 57.406 39.304 57.454 ;
        RECT 22.29 57.452 39.258 57.5 ;
        RECT 22.244 57.498 39.212 57.546 ;
        RECT 22.198 57.544 39.166 57.592 ;
        RECT 22.152 57.59 39.12 57.638 ;
        RECT 22.106 57.636 39.074 57.684 ;
        RECT 22.06 57.682 39.028 57.73 ;
        RECT 22.014 57.728 38.982 57.776 ;
        RECT 21.968 57.774 38.936 57.822 ;
        RECT 21.922 57.82 38.89 57.868 ;
        RECT 21.876 57.866 38.844 57.914 ;
        RECT 21.83 57.912 38.798 57.96 ;
        RECT 21.784 57.958 38.752 58.006 ;
        RECT 21.738 58.004 38.706 58.052 ;
        RECT 21.692 58.05 38.66 58.098 ;
        RECT 21.646 58.096 38.614 58.144 ;
        RECT 21.6 58.142 38.568 58.19 ;
        RECT 21.554 58.188 38.522 58.236 ;
        RECT 21.508 58.234 38.476 58.282 ;
        RECT 21.462 58.28 38.43 58.328 ;
        RECT 21.416 58.326 38.384 58.374 ;
        RECT 21.37 58.372 38.338 58.42 ;
        RECT 21.324 58.418 38.292 58.466 ;
        RECT 21.278 58.464 38.246 58.512 ;
        RECT 21.232 58.51 38.2 58.558 ;
        RECT 21.186 58.556 38.154 58.604 ;
        RECT 21.14 58.602 38.108 58.65 ;
        RECT 21.094 58.648 38.062 58.696 ;
        RECT 21.048 58.694 38.016 58.742 ;
        RECT 21.002 58.74 37.97 58.788 ;
        RECT 20.956 58.786 37.924 58.834 ;
        RECT 20.91 58.832 37.878 58.88 ;
        RECT 20.864 58.878 37.832 58.926 ;
        RECT 20.818 58.924 37.786 58.972 ;
        RECT 20.772 58.97 37.74 59.018 ;
        RECT 20.726 59.016 37.694 59.064 ;
        RECT 20.68 59.062 37.648 59.11 ;
        RECT 20.634 59.108 37.602 59.156 ;
        RECT 20.588 59.154 37.556 59.202 ;
        RECT 20.542 59.2 37.51 59.248 ;
        RECT 20.496 59.246 37.464 59.294 ;
        RECT 20.45 59.292 37.418 59.34 ;
        RECT 20.404 59.338 37.372 59.386 ;
        RECT 20.358 59.384 37.326 59.432 ;
        RECT 20.312 59.43 37.28 59.478 ;
        RECT 20.266 59.476 37.234 59.524 ;
        RECT 20.22 59.522 37.188 59.57 ;
        RECT 20.174 59.568 37.142 59.616 ;
        RECT 20.128 59.614 37.096 59.662 ;
        RECT 20.082 59.66 37.05 59.708 ;
        RECT 20.036 59.706 37.004 59.754 ;
        RECT 19.99 59.752 36.958 59.8 ;
        RECT 19.944 59.798 36.912 59.846 ;
        RECT 19.898 59.844 36.866 59.892 ;
        RECT 19.852 59.89 36.82 59.938 ;
        RECT 19.806 59.936 36.774 59.984 ;
        RECT 19.76 59.982 36.728 60.03 ;
        RECT 19.714 60.028 36.682 60.076 ;
        RECT 19.668 60.074 36.636 60.122 ;
        RECT 19.622 60.12 36.59 60.168 ;
        RECT 19.576 60.166 36.544 60.214 ;
        RECT 19.53 60.212 36.498 60.26 ;
        RECT 19.484 60.258 36.452 60.306 ;
        RECT 19.438 60.304 36.406 60.352 ;
        RECT 19.392 60.35 36.36 60.398 ;
        RECT 19.346 60.396 36.314 60.444 ;
        RECT 19.3 60.442 36.268 60.49 ;
        RECT 19.254 60.488 36.222 60.536 ;
        RECT 19.208 60.534 36.176 60.582 ;
        RECT 19.162 60.58 36.13 60.628 ;
        RECT 19.116 60.626 36.084 60.674 ;
        RECT 19.07 60.672 36.038 60.72 ;
        RECT 19.024 60.718 35.992 60.766 ;
        RECT 18.978 60.764 35.946 60.812 ;
        RECT 18.932 60.81 35.9 60.858 ;
        RECT 18.886 60.856 35.854 60.904 ;
        RECT 18.84 60.902 35.808 60.95 ;
        RECT 18.794 60.948 35.762 60.996 ;
        RECT 18.748 60.994 35.716 61.042 ;
        RECT 18.702 61.04 35.67 61.088 ;
        RECT 18.656 61.086 35.624 61.134 ;
        RECT 18.61 61.132 35.578 61.18 ;
        RECT 18.564 61.178 35.532 61.226 ;
        RECT 18.518 61.224 35.486 61.272 ;
        RECT 18.472 61.27 35.44 61.318 ;
        RECT 18.426 61.316 35.394 61.364 ;
        RECT 18.38 61.362 35.348 61.41 ;
        RECT 18.334 61.408 35.302 61.456 ;
        RECT 18.288 61.454 35.256 61.502 ;
        RECT 18.242 61.5 35.21 61.548 ;
        RECT 18.196 61.546 35.164 61.594 ;
        RECT 18.15 61.592 35.118 61.64 ;
        RECT 18.104 61.638 35.072 61.686 ;
        RECT 18.058 61.684 35.026 61.732 ;
        RECT 18.012 61.73 34.98 61.778 ;
        RECT 17.966 61.776 34.934 61.824 ;
        RECT 17.92 61.822 34.888 61.87 ;
        RECT 17.874 61.868 34.842 61.916 ;
        RECT 17.828 61.914 34.796 61.962 ;
        RECT 17.782 61.96 34.75 62.008 ;
        RECT 17.736 62.006 34.704 62.054 ;
        RECT 17.69 62.052 34.658 62.1 ;
        RECT 17.644 62.098 34.612 62.146 ;
        RECT 17.598 62.144 34.566 62.192 ;
        RECT 17.552 62.19 34.52 62.238 ;
        RECT 17.506 62.236 34.474 62.284 ;
        RECT 17.46 62.282 34.428 62.33 ;
        RECT 17.414 62.328 34.382 62.376 ;
        RECT 17.368 62.374 34.336 62.422 ;
        RECT 17.322 62.42 34.29 62.468 ;
        RECT 17.276 62.466 34.244 62.514 ;
        RECT 17.23 62.512 34.198 62.56 ;
        RECT 17.184 62.558 34.152 62.606 ;
        RECT 17.138 62.604 34.106 62.652 ;
        RECT 17.092 62.65 34.06 62.698 ;
        RECT 17.046 62.696 34.014 62.744 ;
        RECT 17 62.742 33.968 62.79 ;
        RECT 17 62.742 33.922 62.836 ;
        RECT 17 62.742 33.876 62.882 ;
        RECT 17 62.742 33.83 62.928 ;
        RECT 17 62.742 33.784 62.974 ;
        RECT 17 62.742 33.738 63.02 ;
        RECT 17 62.742 33.692 63.066 ;
        RECT 17 62.742 33.646 63.112 ;
        RECT 17 62.742 33.6 63.158 ;
        RECT 17 62.742 33.554 63.204 ;
        RECT 17 62.742 33.508 63.25 ;
        RECT 17 62.742 33.462 63.296 ;
        RECT 17 62.742 33.416 63.342 ;
        RECT 17 62.742 33.37 63.388 ;
        RECT 17 62.742 33.324 63.434 ;
        RECT 17 62.742 33.278 63.48 ;
        RECT 17 62.742 33.232 63.526 ;
        RECT 17 62.742 33.186 63.572 ;
        RECT 17 62.742 33.14 63.618 ;
        RECT 17 62.742 33.094 63.664 ;
        RECT 17 62.742 33.048 63.71 ;
        RECT 17 62.742 33.002 63.756 ;
        RECT 17 62.742 32.956 63.802 ;
        RECT 17 62.742 32.91 63.848 ;
        RECT 17 62.742 32.864 63.894 ;
        RECT 17 62.742 32.818 63.94 ;
        RECT 17 62.742 32.772 63.986 ;
        RECT 17 62.742 32.726 64.032 ;
        RECT 17 62.742 32.68 64.078 ;
        RECT 17 62.742 32.634 64.124 ;
        RECT 17 62.742 32.588 64.17 ;
        RECT 17 62.742 32.542 64.216 ;
        RECT 17 62.742 32.496 64.262 ;
        RECT 17 62.742 32.45 64.308 ;
        RECT 17 62.742 32.404 64.354 ;
        RECT 17 62.742 32.358 64.4 ;
        RECT 17 62.742 32.312 64.446 ;
        RECT 17 62.742 32.266 64.492 ;
        RECT 17 62.742 32.22 64.538 ;
        RECT 17 62.742 32.174 64.584 ;
        RECT 17 62.742 32.128 64.63 ;
        RECT 17 62.742 32.082 64.676 ;
        RECT 17 62.742 32.036 64.722 ;
        RECT 17 62.742 31.99 64.768 ;
        RECT 17 62.742 31.944 64.814 ;
        RECT 17 62.742 31.898 64.86 ;
        RECT 17 62.742 31.852 64.906 ;
        RECT 17 62.742 31.806 64.952 ;
        RECT 17 62.742 31.76 64.998 ;
        RECT 17 62.742 31.714 65.044 ;
        RECT 17 62.742 31.668 65.09 ;
        RECT 17 62.742 31.622 65.136 ;
        RECT 17 62.742 31.576 65.182 ;
        RECT 17 62.742 31.53 65.228 ;
        RECT 17 62.742 31.484 65.274 ;
        RECT 17 62.742 31.438 65.32 ;
        RECT 17 62.742 31.392 65.366 ;
        RECT 17 62.742 31.346 65.412 ;
        RECT 17 62.742 31.3 65.458 ;
        RECT 17 62.742 31.254 65.504 ;
        RECT 17 62.742 31.208 65.55 ;
        RECT 17 62.742 31.162 65.596 ;
        RECT 17 62.742 31.116 65.642 ;
        RECT 17 62.742 31.07 65.688 ;
        RECT 17 62.742 31.024 65.734 ;
        RECT 17 62.742 30.978 65.78 ;
        RECT 17 62.742 30.932 65.826 ;
        RECT 17 62.742 30.886 65.872 ;
        RECT 17 62.742 30.84 65.918 ;
        RECT 17 62.742 30.794 65.964 ;
        RECT 17 62.742 30.748 66.01 ;
        RECT 17 62.742 30.702 66.056 ;
        RECT 17 62.742 30.656 66.102 ;
        RECT 17 62.742 30.61 66.148 ;
        RECT 17 62.742 30.564 66.194 ;
        RECT 17 62.742 30.518 66.24 ;
        RECT 17 62.742 30.472 66.286 ;
        RECT 17 62.742 30.426 66.332 ;
        RECT 17 62.742 30.38 66.378 ;
        RECT 17 62.742 30.334 66.424 ;
        RECT 17 62.742 30.288 66.47 ;
        RECT 17 62.742 30.242 66.516 ;
        RECT 17 62.742 30.196 66.562 ;
        RECT 17 62.742 30.15 66.608 ;
        RECT 17 62.742 30.104 66.654 ;
        RECT 17 62.742 30.058 66.7 ;
        RECT 17 62.742 30.012 66.746 ;
        RECT 17 62.742 29.966 66.792 ;
        RECT 17 62.742 29.92 66.838 ;
        RECT 17 62.742 29.874 66.884 ;
        RECT 17 62.742 29.828 66.93 ;
        RECT 17 62.742 29.782 66.976 ;
        RECT 17 62.742 29.736 67.022 ;
        RECT 17 62.742 29.69 67.068 ;
        RECT 17 62.742 29.644 67.114 ;
        RECT 17 62.742 29.598 67.16 ;
        RECT 17 62.742 29.552 67.206 ;
        RECT 17 62.742 29.506 67.252 ;
        RECT 17 62.742 29.46 67.298 ;
        RECT 17 62.742 29.414 67.344 ;
        RECT 17 62.742 29.368 67.39 ;
        RECT 17 62.742 29.322 67.436 ;
        RECT 17 62.742 29.276 67.482 ;
        RECT 17 62.742 29.23 67.528 ;
        RECT 17 62.742 29.184 67.574 ;
        RECT 17 62.742 29.138 67.62 ;
        RECT 17 62.742 29.092 67.666 ;
        RECT 17 62.742 29.046 67.712 ;
        RECT 17 62.742 29 110 ;
        RECT 92.47 78.5 110 89.5 ;
        RECT 81.444 89.503 97.024 89.529 ;
        RECT 78.5 92.447 94.034 92.519 ;
        RECT 78.5 92.447 93.988 92.565 ;
        RECT 78.5 92.447 93.942 92.611 ;
        RECT 78.5 92.447 93.896 92.657 ;
        RECT 78.5 92.447 93.85 92.703 ;
        RECT 78.5 92.447 93.804 92.749 ;
        RECT 78.5 92.447 93.758 92.795 ;
        RECT 78.5 92.447 93.712 92.841 ;
        RECT 78.5 92.447 93.666 92.887 ;
        RECT 78.5 92.447 93.62 92.933 ;
        RECT 78.5 92.447 93.574 92.979 ;
        RECT 78.5 92.447 93.528 93.025 ;
        RECT 78.5 92.447 93.482 93.071 ;
        RECT 78.5 92.447 93.436 93.117 ;
        RECT 78.5 92.447 93.39 93.163 ;
        RECT 78.5 92.447 93.344 93.209 ;
        RECT 78.5 92.447 93.298 93.255 ;
        RECT 78.5 92.447 93.252 93.301 ;
        RECT 78.5 92.447 93.206 93.347 ;
        RECT 78.5 92.447 93.16 93.393 ;
        RECT 78.5 92.447 93.114 93.439 ;
        RECT 78.5 92.447 93.068 93.485 ;
        RECT 78.5 92.447 93.022 93.531 ;
        RECT 78.5 92.447 92.976 93.577 ;
        RECT 78.5 92.447 92.93 93.623 ;
        RECT 78.5 92.447 92.884 93.669 ;
        RECT 78.5 92.447 92.838 93.715 ;
        RECT 78.5 92.447 92.792 93.761 ;
        RECT 78.5 92.447 92.746 93.807 ;
        RECT 78.5 92.447 92.7 93.853 ;
        RECT 78.5 92.447 92.654 93.899 ;
        RECT 78.5 92.447 92.608 93.945 ;
        RECT 78.5 92.447 92.562 93.991 ;
        RECT 78.5 92.447 92.516 94.037 ;
        RECT 78.546 92.401 94.08 92.473 ;
        RECT 92.444 78.513 92.47 94.073 ;
        RECT 78.592 92.355 94.126 92.427 ;
        RECT 92.398 78.549 92.444 94.109 ;
        RECT 78.638 92.309 94.172 92.381 ;
        RECT 92.352 78.595 92.398 94.155 ;
        RECT 78.684 92.263 94.218 92.335 ;
        RECT 92.306 78.641 92.352 94.201 ;
        RECT 78.73 92.217 94.264 92.289 ;
        RECT 92.26 78.687 92.306 94.247 ;
        RECT 78.776 92.171 94.31 92.243 ;
        RECT 92.214 78.733 92.26 94.293 ;
        RECT 78.822 92.125 94.356 92.197 ;
        RECT 92.168 78.779 92.214 94.339 ;
        RECT 78.868 92.079 94.402 92.151 ;
        RECT 92.122 78.825 92.168 94.385 ;
        RECT 78.914 92.033 94.448 92.105 ;
        RECT 92.076 78.871 92.122 94.431 ;
        RECT 78.96 91.987 94.494 92.059 ;
        RECT 92.03 78.917 92.076 94.477 ;
        RECT 79.006 91.941 94.54 92.013 ;
        RECT 91.984 78.963 92.03 94.523 ;
        RECT 79.052 91.895 94.586 91.967 ;
        RECT 91.938 79.009 91.984 94.569 ;
        RECT 79.098 91.849 94.632 91.921 ;
        RECT 91.892 79.055 91.938 94.615 ;
        RECT 79.144 91.803 94.678 91.875 ;
        RECT 91.846 79.101 91.892 94.661 ;
        RECT 79.19 91.757 94.724 91.829 ;
        RECT 91.8 79.147 91.846 94.707 ;
        RECT 79.236 91.711 94.77 91.783 ;
        RECT 91.754 79.193 91.8 94.753 ;
        RECT 79.282 91.665 94.816 91.737 ;
        RECT 91.708 79.239 91.754 94.799 ;
        RECT 79.328 91.619 94.862 91.691 ;
        RECT 91.662 79.285 91.708 94.845 ;
        RECT 79.374 91.573 94.908 91.645 ;
        RECT 91.616 79.331 91.662 94.891 ;
        RECT 79.42 91.527 94.954 91.599 ;
        RECT 91.57 79.377 91.616 94.937 ;
        RECT 79.466 91.481 95 91.553 ;
        RECT 91.524 79.423 91.57 94.983 ;
        RECT 79.512 91.435 95.046 91.507 ;
        RECT 91.478 79.469 91.524 95.029 ;
        RECT 79.558 91.389 95.092 91.461 ;
        RECT 91.432 79.515 91.478 95.075 ;
        RECT 79.604 91.343 95.138 91.415 ;
        RECT 91.386 79.561 91.432 95.121 ;
        RECT 79.65 91.297 95.184 91.369 ;
        RECT 91.34 79.607 91.386 95.167 ;
        RECT 79.696 91.251 95.23 91.323 ;
        RECT 91.294 79.653 91.34 95.213 ;
        RECT 79.742 91.205 95.276 91.277 ;
        RECT 91.248 79.699 91.294 95.259 ;
        RECT 79.788 91.159 95.322 91.231 ;
        RECT 91.202 79.745 91.248 95.305 ;
        RECT 79.834 91.113 95.368 91.185 ;
        RECT 91.156 79.791 91.202 95.351 ;
        RECT 79.88 91.067 95.414 91.139 ;
        RECT 91.11 79.837 91.156 95.397 ;
        RECT 79.926 91.021 95.46 91.093 ;
        RECT 91.064 79.883 91.11 95.443 ;
        RECT 79.972 90.975 95.506 91.047 ;
        RECT 91.018 79.929 91.064 95.489 ;
        RECT 80.018 90.929 95.552 91.001 ;
        RECT 90.972 79.975 91.018 95.535 ;
        RECT 80.064 90.883 95.598 90.955 ;
        RECT 90.926 80.021 90.972 95.581 ;
        RECT 80.11 90.837 95.644 90.909 ;
        RECT 90.88 80.067 90.926 95.627 ;
        RECT 80.156 90.791 95.69 90.863 ;
        RECT 90.834 80.113 90.88 95.673 ;
        RECT 80.202 90.745 95.736 90.817 ;
        RECT 90.788 80.159 90.834 95.719 ;
        RECT 80.248 90.699 95.782 90.771 ;
        RECT 90.742 80.205 90.788 95.765 ;
        RECT 80.294 90.653 95.828 90.725 ;
        RECT 90.696 80.251 90.742 95.811 ;
        RECT 80.34 90.607 95.874 90.679 ;
        RECT 90.65 80.297 90.696 95.857 ;
        RECT 80.386 90.561 95.92 90.633 ;
        RECT 90.604 80.343 90.65 95.903 ;
        RECT 80.432 90.515 95.966 90.587 ;
        RECT 90.558 80.389 90.604 95.949 ;
        RECT 80.478 90.469 96.012 90.541 ;
        RECT 90.512 80.435 90.558 95.995 ;
        RECT 80.524 90.423 96.058 90.495 ;
        RECT 90.466 80.481 90.512 96.041 ;
        RECT 80.57 90.377 96.104 90.449 ;
        RECT 90.42 80.527 90.466 96.087 ;
        RECT 80.616 90.331 96.15 90.403 ;
        RECT 90.374 80.573 90.42 96.133 ;
        RECT 80.662 90.285 96.196 90.357 ;
        RECT 90.328 80.619 90.374 96.179 ;
        RECT 80.708 90.239 96.242 90.311 ;
        RECT 90.282 80.665 90.328 96.225 ;
        RECT 80.754 90.193 96.288 90.265 ;
        RECT 90.236 80.711 90.282 96.271 ;
        RECT 80.8 90.147 96.334 90.219 ;
        RECT 90.19 80.757 90.236 96.317 ;
        RECT 80.846 90.101 96.38 90.173 ;
        RECT 90.144 80.803 90.19 96.363 ;
        RECT 80.892 90.055 96.426 90.127 ;
        RECT 90.098 80.849 90.144 96.409 ;
        RECT 80.938 90.009 96.472 90.081 ;
        RECT 90.052 80.895 90.098 96.455 ;
        RECT 80.984 89.963 96.518 90.035 ;
        RECT 90.006 80.941 90.052 96.501 ;
        RECT 81.03 89.917 96.564 89.989 ;
        RECT 89.96 80.987 90.006 96.547 ;
        RECT 81.076 89.871 96.61 89.943 ;
        RECT 89.914 81.033 89.96 96.593 ;
        RECT 81.122 89.825 96.656 89.897 ;
        RECT 89.868 81.079 89.914 96.639 ;
        RECT 81.168 89.779 96.702 89.851 ;
        RECT 89.822 81.125 89.868 96.685 ;
        RECT 81.214 89.733 96.748 89.805 ;
        RECT 89.776 81.171 89.822 96.731 ;
        RECT 81.26 89.687 96.794 89.759 ;
        RECT 89.73 81.217 89.776 96.777 ;
        RECT 81.306 89.641 96.84 89.713 ;
        RECT 89.684 81.263 89.73 96.823 ;
        RECT 81.352 89.595 96.886 89.667 ;
        RECT 89.638 81.309 89.684 96.869 ;
        RECT 81.398 89.549 96.932 89.621 ;
        RECT 89.592 81.355 89.638 96.915 ;
        RECT 81.444 89.503 96.978 89.575 ;
        RECT 89.546 81.401 89.592 96.961 ;
        RECT 81.49 89.457 97.03 89.503 ;
        RECT 89.5 81.447 89.546 97.007 ;
        RECT 78.5 92.447 89.5 110 ;
        RECT 81.536 89.411 110 89.5 ;
        RECT 89.494 81.473 89.5 110 ;
        RECT 81.582 89.365 110 89.5 ;
        RECT 89.448 81.499 89.5 110 ;
        RECT 81.628 89.319 110 89.5 ;
        RECT 89.402 81.545 89.5 110 ;
        RECT 81.674 89.273 110 89.5 ;
        RECT 89.356 81.591 89.5 110 ;
        RECT 81.72 89.227 110 89.5 ;
        RECT 89.31 81.637 89.5 110 ;
        RECT 81.766 89.181 110 89.5 ;
        RECT 89.264 81.683 89.5 110 ;
        RECT 81.812 89.135 110 89.5 ;
        RECT 89.218 81.729 89.5 110 ;
        RECT 81.858 89.089 110 89.5 ;
        RECT 89.172 81.775 89.5 110 ;
        RECT 81.904 89.043 110 89.5 ;
        RECT 89.126 81.821 89.5 110 ;
        RECT 81.95 88.997 110 89.5 ;
        RECT 89.08 81.867 89.5 110 ;
        RECT 81.996 88.951 110 89.5 ;
        RECT 89.034 81.913 89.5 110 ;
        RECT 82.042 88.905 110 89.5 ;
        RECT 88.988 81.959 89.5 110 ;
        RECT 82.088 88.859 110 89.5 ;
        RECT 88.942 82.005 89.5 110 ;
        RECT 82.134 88.813 110 89.5 ;
        RECT 88.896 82.051 89.5 110 ;
        RECT 82.18 88.767 110 89.5 ;
        RECT 88.85 82.097 89.5 110 ;
        RECT 82.226 88.721 110 89.5 ;
        RECT 88.804 82.143 89.5 110 ;
        RECT 82.272 88.675 110 89.5 ;
        RECT 88.758 82.189 89.5 110 ;
        RECT 82.318 88.629 110 89.5 ;
        RECT 88.712 82.235 89.5 110 ;
        RECT 82.364 88.583 110 89.5 ;
        RECT 88.666 82.281 89.5 110 ;
        RECT 82.41 88.537 110 89.5 ;
        RECT 88.62 82.327 89.5 110 ;
        RECT 82.456 88.491 110 89.5 ;
        RECT 88.574 82.373 89.5 110 ;
        RECT 82.502 88.445 110 89.5 ;
        RECT 88.528 82.419 89.5 110 ;
        RECT 82.548 88.399 110 89.5 ;
        RECT 88.482 82.465 89.5 110 ;
        RECT 82.594 88.353 110 89.5 ;
        RECT 88.436 82.511 89.5 110 ;
        RECT 82.64 88.307 110 89.5 ;
        RECT 88.39 82.557 89.5 110 ;
        RECT 82.686 88.261 110 89.5 ;
        RECT 88.344 82.603 89.5 110 ;
        RECT 82.732 88.215 110 89.5 ;
        RECT 88.298 82.649 89.5 110 ;
        RECT 82.778 88.169 110 89.5 ;
        RECT 88.252 82.695 89.5 110 ;
        RECT 82.824 88.123 110 89.5 ;
        RECT 88.206 82.741 89.5 110 ;
        RECT 82.87 88.077 110 89.5 ;
        RECT 88.16 82.787 89.5 110 ;
        RECT 82.916 88.031 110 89.5 ;
        RECT 88.114 82.833 89.5 110 ;
        RECT 82.962 87.985 110 89.5 ;
        RECT 88.068 82.879 89.5 110 ;
        RECT 83.008 87.939 110 89.5 ;
        RECT 88.022 82.925 89.5 110 ;
        RECT 83.054 87.893 110 89.5 ;
        RECT 87.976 82.971 89.5 110 ;
        RECT 83.1 87.847 110 89.5 ;
        RECT 87.93 83.017 89.5 110 ;
        RECT 83.146 87.801 110 89.5 ;
        RECT 87.884 83.063 89.5 110 ;
        RECT 83.192 87.755 110 89.5 ;
        RECT 87.838 83.109 89.5 110 ;
        RECT 83.238 87.709 110 89.5 ;
        RECT 87.792 83.155 89.5 110 ;
        RECT 83.284 87.663 110 89.5 ;
        RECT 87.746 83.201 89.5 110 ;
        RECT 83.33 87.617 110 89.5 ;
        RECT 87.7 83.247 89.5 110 ;
        RECT 83.376 87.571 110 89.5 ;
        RECT 87.654 83.293 89.5 110 ;
        RECT 83.422 87.525 110 89.5 ;
        RECT 87.608 83.339 89.5 110 ;
        RECT 83.468 87.479 110 89.5 ;
        RECT 87.562 83.385 89.5 110 ;
        RECT 83.514 87.433 110 89.5 ;
        RECT 87.516 83.431 89.5 110 ;
        RECT 83.56 87.387 110 89.5 ;
        RECT 87.47 83.477 89.5 110 ;
        RECT 83.606 87.341 110 89.5 ;
        RECT 87.424 83.523 89.5 110 ;
        RECT 83.652 87.295 110 89.5 ;
        RECT 87.378 83.569 89.5 110 ;
        RECT 83.698 87.249 110 89.5 ;
        RECT 87.332 83.615 89.5 110 ;
        RECT 83.744 87.203 110 89.5 ;
        RECT 87.286 83.661 89.5 110 ;
        RECT 83.79 87.157 110 89.5 ;
        RECT 87.24 83.707 89.5 110 ;
        RECT 83.836 87.111 110 89.5 ;
        RECT 87.194 83.753 89.5 110 ;
        RECT 83.882 87.065 110 89.5 ;
        RECT 87.148 83.799 89.5 110 ;
        RECT 83.928 87.019 110 89.5 ;
        RECT 87.102 83.845 89.5 110 ;
        RECT 83.974 86.973 110 89.5 ;
        RECT 87.056 83.891 89.5 110 ;
        RECT 84.02 86.927 110 89.5 ;
        RECT 87.01 83.937 89.5 110 ;
        RECT 84.066 86.881 110 89.5 ;
        RECT 86.964 83.983 89.5 110 ;
        RECT 84.112 86.835 110 89.5 ;
        RECT 86.918 84.029 89.5 110 ;
        RECT 84.158 86.789 110 89.5 ;
        RECT 86.872 84.075 89.5 110 ;
        RECT 84.204 86.743 110 89.5 ;
        RECT 86.826 84.121 89.5 110 ;
        RECT 84.25 86.697 110 89.5 ;
        RECT 86.78 84.167 89.5 110 ;
        RECT 84.296 86.651 110 89.5 ;
        RECT 86.734 84.213 89.5 110 ;
        RECT 84.342 86.605 110 89.5 ;
        RECT 86.688 84.259 89.5 110 ;
        RECT 84.388 86.559 110 89.5 ;
        RECT 86.642 84.305 89.5 110 ;
        RECT 84.434 86.513 110 89.5 ;
        RECT 86.596 84.351 89.5 110 ;
        RECT 84.48 86.467 110 89.5 ;
        RECT 86.55 84.397 89.5 110 ;
        RECT 84.526 86.421 110 89.5 ;
        RECT 86.504 84.443 89.5 110 ;
        RECT 84.572 86.375 110 89.5 ;
        RECT 86.458 84.489 89.5 110 ;
        RECT 84.618 86.329 110 89.5 ;
        RECT 86.412 84.535 89.5 110 ;
        RECT 84.664 86.283 110 89.5 ;
        RECT 86.366 84.581 89.5 110 ;
        RECT 84.71 86.237 110 89.5 ;
        RECT 86.32 84.627 89.5 110 ;
        RECT 84.756 86.191 110 89.5 ;
        RECT 86.274 84.673 89.5 110 ;
        RECT 84.802 86.145 110 89.5 ;
        RECT 86.228 84.719 89.5 110 ;
        RECT 84.848 86.099 110 89.5 ;
        RECT 86.182 84.765 89.5 110 ;
        RECT 84.894 86.053 110 89.5 ;
        RECT 86.136 84.811 89.5 110 ;
        RECT 84.94 86.007 110 89.5 ;
        RECT 86.09 84.857 89.5 110 ;
        RECT 84.986 85.961 110 89.5 ;
        RECT 86.044 84.903 89.5 110 ;
        RECT 85.032 85.915 110 89.5 ;
        RECT 85.998 84.949 89.5 110 ;
        RECT 85.078 85.869 110 89.5 ;
        RECT 85.952 84.995 89.5 110 ;
        RECT 85.124 85.823 110 89.5 ;
        RECT 85.906 85.041 89.5 110 ;
        RECT 85.17 85.777 110 89.5 ;
        RECT 85.86 85.087 89.5 110 ;
        RECT 85.216 85.731 110 89.5 ;
        RECT 85.814 85.133 89.5 110 ;
        RECT 85.262 85.685 110 89.5 ;
        RECT 85.768 85.179 89.5 110 ;
        RECT 85.308 85.639 110 89.5 ;
        RECT 85.722 85.225 89.5 110 ;
        RECT 85.354 85.593 110 89.5 ;
        RECT 85.676 85.271 89.5 110 ;
        RECT 85.4 85.547 110 89.5 ;
        RECT 85.63 85.317 89.5 110 ;
        RECT 85.446 85.501 110 89.5 ;
        RECT 85.584 85.363 89.5 110 ;
        RECT 85.492 85.455 110 89.5 ;
        RECT 85.538 85.409 89.5 110 ;
        RECT 10.032 49.46 27 49.508 ;
        RECT 9.986 49.506 26.954 49.554 ;
        RECT 9.94 49.552 26.908 49.6 ;
        RECT 9.894 49.598 26.862 49.646 ;
        RECT 9.848 49.644 26.816 49.692 ;
        RECT 9.802 49.69 26.77 49.738 ;
        RECT 9.756 49.736 26.724 49.784 ;
        RECT 9.71 49.782 26.678 49.83 ;
        RECT 9.664 49.828 26.632 49.876 ;
        RECT 9.618 49.874 26.586 49.922 ;
        RECT 9.572 49.92 26.54 49.968 ;
        RECT 9.526 49.966 26.494 50.014 ;
        RECT 9.48 50.012 26.448 50.06 ;
        RECT 9.434 50.058 26.402 50.106 ;
        RECT 9.388 50.104 26.356 50.152 ;
        RECT 9.342 50.15 26.31 50.198 ;
        RECT 9.296 50.196 26.264 50.244 ;
        RECT 9.25 50.242 26.218 50.29 ;
        RECT 9.204 50.288 26.172 50.336 ;
        RECT 9.158 50.334 26.126 50.382 ;
        RECT 9.112 50.38 26.08 50.428 ;
        RECT 9.066 50.426 26.034 50.474 ;
        RECT 9.02 50.472 25.988 50.52 ;
        RECT 8.974 50.518 25.942 50.566 ;
        RECT 8.928 50.564 25.896 50.612 ;
        RECT 8.882 50.61 25.85 50.658 ;
        RECT 8.836 50.656 25.804 50.704 ;
        RECT 8.79 50.702 25.758 50.75 ;
        RECT 8.744 50.748 25.712 50.796 ;
        RECT 8.698 50.794 25.666 50.842 ;
        RECT 8.652 50.84 25.62 50.888 ;
        RECT 8.606 50.886 25.574 50.934 ;
        RECT 8.56 50.932 25.528 50.98 ;
        RECT 8.514 50.978 25.482 51.026 ;
        RECT 8.468 51.024 25.436 51.072 ;
        RECT 8.422 51.07 25.39 51.118 ;
        RECT 8.376 51.116 25.344 51.164 ;
        RECT 8.33 51.162 25.298 51.21 ;
        RECT 8.284 51.208 25.252 51.256 ;
        RECT 8.238 51.254 25.206 51.302 ;
        RECT 8.192 51.3 25.16 51.348 ;
        RECT 8.146 51.346 25.114 51.394 ;
        RECT 8.1 51.392 25.068 51.44 ;
        RECT 8.054 51.438 25.022 51.486 ;
        RECT 8.008 51.484 24.976 51.532 ;
        RECT 7.962 51.53 24.93 51.578 ;
        RECT 7.916 51.576 24.884 51.624 ;
        RECT 7.87 51.622 24.838 51.67 ;
        RECT 7.824 51.668 24.792 51.716 ;
        RECT 7.778 51.714 24.746 51.762 ;
        RECT 7.732 51.76 24.7 51.808 ;
        RECT 7.686 51.806 24.654 51.854 ;
        RECT 7.64 51.852 24.608 51.9 ;
        RECT 7.594 51.898 24.562 51.946 ;
        RECT 7.548 51.944 24.516 51.992 ;
        RECT 7.502 51.99 24.47 52.038 ;
        RECT 7.456 52.036 24.424 52.084 ;
        RECT 7.41 52.082 24.378 52.13 ;
        RECT 7.364 52.128 24.332 52.176 ;
        RECT 7.318 52.174 24.286 52.222 ;
        RECT 7.272 52.22 24.24 52.268 ;
        RECT 7.226 52.266 24.194 52.314 ;
        RECT 7.18 52.312 24.148 52.36 ;
        RECT 7.134 52.358 24.102 52.406 ;
        RECT 7.088 52.404 24.056 52.452 ;
        RECT 7.042 52.45 24.01 52.498 ;
        RECT 6.996 52.496 23.964 52.544 ;
        RECT 6.95 52.542 23.918 52.59 ;
        RECT 6.904 52.588 23.872 52.636 ;
        RECT 6.858 52.634 23.826 52.682 ;
        RECT 6.812 52.68 23.78 52.728 ;
        RECT 6.766 52.726 23.734 52.774 ;
        RECT 6.72 52.772 23.688 52.82 ;
        RECT 6.674 52.818 23.642 52.866 ;
        RECT 6.628 52.864 23.596 52.912 ;
        RECT 6.582 52.91 23.55 52.958 ;
        RECT 6.536 52.956 23.504 53.004 ;
        RECT 6.49 53.002 23.458 53.05 ;
        RECT 6.444 53.048 23.412 53.096 ;
        RECT 6.398 53.094 23.366 53.142 ;
        RECT 6.352 53.14 23.32 53.188 ;
        RECT 6.306 53.186 23.274 53.234 ;
        RECT 6.26 53.232 23.228 53.28 ;
        RECT 6.214 53.278 23.182 53.326 ;
        RECT 6.168 53.324 23.136 53.372 ;
        RECT 6.122 53.37 23.09 53.418 ;
        RECT 6.076 53.416 23.044 53.464 ;
        RECT 6.03 53.462 22.998 53.51 ;
        RECT 5.984 53.508 22.952 53.556 ;
        RECT 5.938 53.554 22.906 53.602 ;
        RECT 5.892 53.6 22.86 53.648 ;
        RECT 5.846 53.646 22.814 53.694 ;
        RECT 5.8 53.692 22.768 53.74 ;
        RECT 5.754 53.738 22.722 53.786 ;
        RECT 5.708 53.784 22.676 53.832 ;
        RECT 5.662 53.83 22.63 53.878 ;
        RECT 5.616 53.876 22.584 53.924 ;
        RECT 5.57 53.922 22.538 53.97 ;
        RECT 5.524 53.968 22.492 54.016 ;
        RECT 5.478 54.014 22.446 54.062 ;
        RECT 5.432 54.06 22.4 54.108 ;
        RECT 5.386 54.106 22.354 54.154 ;
        RECT 5.34 54.152 22.308 54.2 ;
        RECT 5.294 54.198 22.262 54.246 ;
        RECT 5.248 54.244 22.216 54.292 ;
        RECT 5.202 54.29 22.17 54.338 ;
        RECT 5.156 54.336 22.124 54.384 ;
        RECT 5.11 54.382 22.078 54.43 ;
        RECT 5.064 54.428 22.032 54.476 ;
        RECT 5.018 54.474 21.986 54.522 ;
        RECT 4.972 54.52 21.94 54.568 ;
        RECT 4.926 54.566 21.894 54.614 ;
        RECT 4.88 54.612 21.848 54.66 ;
        RECT 4.834 54.658 21.802 54.706 ;
        RECT 4.788 54.704 21.756 54.752 ;
        RECT 4.742 54.75 21.71 54.798 ;
        RECT 4.696 54.796 21.664 54.844 ;
        RECT 4.65 54.842 21.618 54.89 ;
        RECT 4.604 54.888 21.572 54.936 ;
        RECT 4.558 54.934 21.526 54.982 ;
        RECT 4.512 54.98 21.48 55.028 ;
        RECT 4.466 55.026 21.434 55.074 ;
        RECT 4.42 55.072 21.388 55.12 ;
        RECT 4.374 55.118 21.342 55.166 ;
        RECT 4.328 55.164 21.296 55.212 ;
        RECT 4.282 55.21 21.25 55.258 ;
        RECT 4.236 55.256 21.204 55.304 ;
        RECT 4.19 55.302 21.158 55.35 ;
        RECT 4.144 55.348 21.112 55.396 ;
        RECT 4.098 55.394 21.066 55.442 ;
        RECT 4.052 55.44 21.02 55.488 ;
        RECT 4.006 55.486 20.974 55.534 ;
        RECT 3.96 55.532 20.928 55.58 ;
        RECT 3.914 55.578 20.882 55.626 ;
        RECT 3.868 55.624 20.836 55.672 ;
        RECT 3.822 55.67 20.79 55.718 ;
        RECT 3.776 55.716 20.744 55.764 ;
        RECT 3.73 55.762 20.698 55.81 ;
        RECT 3.684 55.808 20.652 55.856 ;
        RECT 3.638 55.854 20.606 55.902 ;
        RECT 3.592 55.9 20.56 55.948 ;
        RECT 3.546 55.946 20.514 55.994 ;
        RECT 3.5 55.992 20.468 56.04 ;
        RECT 3.5 55.992 20.422 56.086 ;
        RECT 3.5 55.992 20.376 56.132 ;
        RECT 3.5 55.992 20.33 56.178 ;
        RECT 3.5 55.992 20.284 56.224 ;
        RECT 3.5 55.992 20.238 56.27 ;
        RECT 3.5 55.992 20.192 56.316 ;
        RECT 3.5 55.992 20.146 56.362 ;
        RECT 3.5 55.992 20.1 56.408 ;
        RECT 3.5 55.992 20.054 56.454 ;
        RECT 3.5 55.992 20.008 56.5 ;
        RECT 3.5 55.992 19.962 56.546 ;
        RECT 3.5 55.992 19.916 56.592 ;
        RECT 3.5 55.992 19.87 56.638 ;
        RECT 3.5 55.992 19.824 56.684 ;
        RECT 3.5 55.992 19.778 56.73 ;
        RECT 3.5 55.992 19.732 56.776 ;
        RECT 3.5 55.992 19.686 56.822 ;
        RECT 3.5 55.992 19.64 56.868 ;
        RECT 3.5 55.992 19.594 56.914 ;
        RECT 3.5 55.992 19.548 56.96 ;
        RECT 3.5 55.992 19.502 57.006 ;
        RECT 3.5 55.992 19.456 57.052 ;
        RECT 3.5 55.992 19.41 57.098 ;
        RECT 3.5 55.992 19.364 57.144 ;
        RECT 3.5 55.992 19.318 57.19 ;
        RECT 3.5 55.992 19.272 57.236 ;
        RECT 3.5 55.992 19.226 57.282 ;
        RECT 3.5 55.992 19.18 57.328 ;
        RECT 3.5 55.992 19.134 57.374 ;
        RECT 3.5 55.992 19.088 57.42 ;
        RECT 3.5 55.992 19.042 57.466 ;
        RECT 3.5 55.992 18.996 57.512 ;
        RECT 3.5 55.992 18.95 57.558 ;
        RECT 3.5 55.992 18.904 57.604 ;
        RECT 3.5 55.992 18.858 57.65 ;
        RECT 3.5 55.992 18.812 57.696 ;
        RECT 3.5 55.992 18.766 57.742 ;
        RECT 3.5 55.992 18.72 57.788 ;
        RECT 3.5 55.992 18.674 57.834 ;
        RECT 3.5 55.992 18.628 57.88 ;
        RECT 3.5 55.992 18.582 57.926 ;
        RECT 3.5 55.992 18.536 57.972 ;
        RECT 3.5 55.992 18.49 58.018 ;
        RECT 3.5 55.992 18.444 58.064 ;
        RECT 3.5 55.992 18.398 58.11 ;
        RECT 3.5 55.992 18.352 58.156 ;
        RECT 3.5 55.992 18.306 58.202 ;
        RECT 3.5 55.992 18.26 58.248 ;
        RECT 3.5 55.992 18.214 58.294 ;
        RECT 3.5 55.992 18.168 58.34 ;
        RECT 3.5 55.992 18.122 58.386 ;
        RECT 3.5 55.992 18.076 58.432 ;
        RECT 3.5 55.992 18.03 58.478 ;
        RECT 3.5 55.992 17.984 58.524 ;
        RECT 3.5 55.992 17.938 58.57 ;
        RECT 3.5 55.992 17.892 58.616 ;
        RECT 3.5 55.992 17.846 58.662 ;
        RECT 3.5 55.992 17.8 58.708 ;
        RECT 3.5 55.992 17.754 58.754 ;
        RECT 3.5 55.992 17.708 58.8 ;
        RECT 3.5 55.992 17.662 58.846 ;
        RECT 3.5 55.992 17.616 58.892 ;
        RECT 3.5 55.992 17.57 58.938 ;
        RECT 3.5 55.992 17.524 58.984 ;
        RECT 3.5 55.992 17.478 59.03 ;
        RECT 3.5 55.992 17.432 59.076 ;
        RECT 3.5 55.992 17.386 59.122 ;
        RECT 3.5 55.992 17.34 59.168 ;
        RECT 3.5 55.992 17.294 59.214 ;
        RECT 3.5 55.992 17.248 59.26 ;
        RECT 3.5 55.992 17.202 59.306 ;
        RECT 3.5 55.992 17.156 59.352 ;
        RECT 3.5 55.992 17.11 59.398 ;
        RECT 3.5 55.992 17.064 59.444 ;
        RECT 3.5 55.992 17.018 59.49 ;
        RECT 3.5 55.992 16.972 59.536 ;
        RECT 3.5 55.992 16.926 59.582 ;
        RECT 3.5 55.992 16.88 59.628 ;
        RECT 3.5 55.992 16.834 59.674 ;
        RECT 3.5 55.992 16.788 59.72 ;
        RECT 3.5 55.992 16.742 59.766 ;
        RECT 3.5 55.992 16.696 59.812 ;
        RECT 3.5 55.992 16.65 59.858 ;
        RECT 3.5 55.992 16.604 59.904 ;
        RECT 3.5 55.992 16.558 59.95 ;
        RECT 3.5 55.992 16.512 59.996 ;
        RECT 3.5 55.992 16.466 60.042 ;
        RECT 3.5 55.992 16.42 60.088 ;
        RECT 3.5 55.992 16.374 60.134 ;
        RECT 3.5 55.992 16.328 60.18 ;
        RECT 3.5 55.992 16.282 60.226 ;
        RECT 3.5 55.992 16.236 60.272 ;
        RECT 3.5 55.992 16.19 60.318 ;
        RECT 3.5 55.992 16.144 60.364 ;
        RECT 3.5 55.992 16.098 60.41 ;
        RECT 3.5 55.992 16.052 60.456 ;
        RECT 3.5 55.992 16.006 60.502 ;
        RECT 3.5 55.992 15.96 60.548 ;
        RECT 3.5 55.992 15.914 60.594 ;
        RECT 3.5 55.992 15.868 60.64 ;
        RECT 3.5 55.992 15.822 60.686 ;
        RECT 3.5 55.992 15.776 60.732 ;
        RECT 3.5 55.992 15.73 60.778 ;
        RECT 3.5 55.992 15.684 60.824 ;
        RECT 3.5 55.992 15.638 60.87 ;
        RECT 3.5 55.992 15.592 60.916 ;
        RECT 3.5 55.992 15.546 60.962 ;
        RECT 3.5 55.992 15.5 110 ;
        RECT 62.764 17 110 29 ;
        RECT 50.758 28.984 67.733 29.024 ;
        RECT 45.836 33.906 62.765 33.971 ;
        RECT 62.718 17.024 62.764 33.994 ;
        RECT 45.79 33.952 62.718 34.04 ;
        RECT 45.882 33.86 62.811 33.947 ;
        RECT 62.672 17.07 62.718 34.04 ;
        RECT 45.744 33.998 62.672 34.086 ;
        RECT 45.928 33.814 62.857 33.901 ;
        RECT 62.626 17.116 62.672 34.086 ;
        RECT 45.698 34.044 62.626 34.132 ;
        RECT 45.974 33.768 62.903 33.855 ;
        RECT 62.58 17.162 62.626 34.132 ;
        RECT 45.652 34.09 62.58 34.178 ;
        RECT 46.02 33.722 62.949 33.809 ;
        RECT 62.534 17.208 62.58 34.178 ;
        RECT 45.606 34.136 62.534 34.224 ;
        RECT 46.066 33.676 62.995 33.763 ;
        RECT 62.488 17.254 62.534 34.224 ;
        RECT 45.56 34.182 62.488 34.27 ;
        RECT 46.112 33.63 63.041 33.717 ;
        RECT 62.442 17.3 62.488 34.27 ;
        RECT 45.514 34.228 62.442 34.316 ;
        RECT 46.158 33.584 63.087 33.671 ;
        RECT 62.396 17.346 62.442 34.316 ;
        RECT 45.468 34.274 62.396 34.362 ;
        RECT 46.204 33.538 63.133 33.625 ;
        RECT 62.35 17.392 62.396 34.362 ;
        RECT 45.422 34.32 62.35 34.408 ;
        RECT 46.25 33.492 63.179 33.579 ;
        RECT 62.304 17.438 62.35 34.408 ;
        RECT 45.376 34.366 62.304 34.454 ;
        RECT 46.296 33.446 63.225 33.533 ;
        RECT 62.258 17.484 62.304 34.454 ;
        RECT 45.33 34.412 62.258 34.5 ;
        RECT 46.342 33.4 63.271 33.487 ;
        RECT 62.212 17.53 62.258 34.5 ;
        RECT 45.284 34.458 62.212 34.546 ;
        RECT 46.388 33.354 63.317 33.441 ;
        RECT 62.166 17.576 62.212 34.546 ;
        RECT 45.238 34.504 62.166 34.592 ;
        RECT 46.434 33.308 63.363 33.395 ;
        RECT 62.12 17.622 62.166 34.592 ;
        RECT 45.192 34.55 62.12 34.638 ;
        RECT 46.48 33.262 63.409 33.349 ;
        RECT 62.074 17.668 62.12 34.638 ;
        RECT 45.146 34.596 62.074 34.684 ;
        RECT 46.526 33.216 63.455 33.303 ;
        RECT 62.028 17.714 62.074 34.684 ;
        RECT 45.1 34.642 62.028 34.73 ;
        RECT 46.572 33.17 63.501 33.257 ;
        RECT 61.982 17.76 62.028 34.73 ;
        RECT 45.054 34.688 61.982 34.776 ;
        RECT 46.618 33.124 63.547 33.211 ;
        RECT 61.936 17.806 61.982 34.776 ;
        RECT 45.008 34.734 61.936 34.822 ;
        RECT 46.664 33.078 63.593 33.165 ;
        RECT 61.89 17.852 61.936 34.822 ;
        RECT 44.962 34.78 61.89 34.868 ;
        RECT 46.71 33.032 63.639 33.119 ;
        RECT 61.844 17.898 61.89 34.868 ;
        RECT 44.916 34.826 61.844 34.914 ;
        RECT 46.756 32.986 63.685 33.073 ;
        RECT 61.798 17.944 61.844 34.914 ;
        RECT 44.87 34.872 61.798 34.96 ;
        RECT 46.802 32.94 63.731 33.027 ;
        RECT 61.752 17.99 61.798 34.96 ;
        RECT 44.824 34.918 61.752 35.006 ;
        RECT 46.848 32.894 63.777 32.981 ;
        RECT 61.706 18.036 61.752 35.006 ;
        RECT 44.778 34.964 61.706 35.052 ;
        RECT 46.894 32.848 63.823 32.935 ;
        RECT 61.66 18.082 61.706 35.052 ;
        RECT 44.732 35.01 61.66 35.098 ;
        RECT 46.94 32.802 63.869 32.889 ;
        RECT 61.614 18.128 61.66 35.098 ;
        RECT 44.686 35.056 61.614 35.144 ;
        RECT 46.986 32.756 63.915 32.843 ;
        RECT 61.568 18.174 61.614 35.144 ;
        RECT 44.64 35.102 61.568 35.19 ;
        RECT 47.032 32.71 63.961 32.797 ;
        RECT 61.522 18.22 61.568 35.19 ;
        RECT 44.594 35.148 61.522 35.236 ;
        RECT 47.078 32.664 64.007 32.751 ;
        RECT 61.476 18.266 61.522 35.236 ;
        RECT 44.548 35.194 61.476 35.282 ;
        RECT 47.124 32.618 64.053 32.705 ;
        RECT 61.43 18.312 61.476 35.282 ;
        RECT 44.502 35.24 61.43 35.328 ;
        RECT 47.17 32.572 64.099 32.659 ;
        RECT 61.384 18.358 61.43 35.328 ;
        RECT 44.456 35.286 61.384 35.374 ;
        RECT 47.216 32.526 64.145 32.613 ;
        RECT 61.338 18.404 61.384 35.374 ;
        RECT 44.41 35.332 61.338 35.42 ;
        RECT 47.262 32.48 64.191 32.567 ;
        RECT 61.292 18.45 61.338 35.42 ;
        RECT 44.364 35.378 61.292 35.466 ;
        RECT 47.308 32.434 64.237 32.521 ;
        RECT 61.246 18.496 61.292 35.466 ;
        RECT 44.318 35.424 61.246 35.512 ;
        RECT 47.354 32.388 64.283 32.475 ;
        RECT 61.2 18.542 61.246 35.512 ;
        RECT 44.272 35.47 61.2 35.558 ;
        RECT 47.4 32.342 64.329 32.429 ;
        RECT 61.154 18.588 61.2 35.558 ;
        RECT 44.226 35.516 61.154 35.604 ;
        RECT 47.446 32.296 64.375 32.383 ;
        RECT 61.108 18.634 61.154 35.604 ;
        RECT 44.18 35.562 61.108 35.65 ;
        RECT 47.492 32.25 64.421 32.337 ;
        RECT 61.062 18.68 61.108 35.65 ;
        RECT 44.134 35.608 61.062 35.696 ;
        RECT 47.538 32.204 64.467 32.291 ;
        RECT 61.016 18.726 61.062 35.696 ;
        RECT 44.088 35.654 61.016 35.742 ;
        RECT 47.584 32.158 64.513 32.245 ;
        RECT 60.97 18.772 61.016 35.742 ;
        RECT 44.042 35.7 60.97 35.788 ;
        RECT 47.63 32.112 64.559 32.199 ;
        RECT 60.924 18.818 60.97 35.788 ;
        RECT 43.996 35.746 60.924 35.834 ;
        RECT 47.676 32.066 64.605 32.153 ;
        RECT 60.878 18.864 60.924 35.834 ;
        RECT 43.95 35.792 60.878 35.88 ;
        RECT 47.722 32.02 64.651 32.107 ;
        RECT 60.832 18.91 60.878 35.88 ;
        RECT 43.904 35.838 60.832 35.926 ;
        RECT 47.768 31.974 64.697 32.061 ;
        RECT 60.786 18.956 60.832 35.926 ;
        RECT 43.858 35.884 60.786 35.972 ;
        RECT 47.814 31.928 64.743 32.015 ;
        RECT 60.74 19.002 60.786 35.972 ;
        RECT 43.812 35.93 60.74 36.018 ;
        RECT 47.86 31.882 64.789 31.969 ;
        RECT 60.694 19.048 60.74 36.018 ;
        RECT 43.766 35.976 60.694 36.064 ;
        RECT 47.906 31.836 64.835 31.923 ;
        RECT 60.648 19.094 60.694 36.064 ;
        RECT 43.72 36.022 60.648 36.11 ;
        RECT 47.952 31.79 64.881 31.877 ;
        RECT 60.602 19.14 60.648 36.11 ;
        RECT 43.674 36.068 60.602 36.156 ;
        RECT 47.998 31.744 64.927 31.831 ;
        RECT 60.556 19.186 60.602 36.156 ;
        RECT 43.628 36.114 60.556 36.202 ;
        RECT 48.044 31.698 64.973 31.785 ;
        RECT 60.51 19.232 60.556 36.202 ;
        RECT 43.582 36.16 60.51 36.248 ;
        RECT 48.09 31.652 65.019 31.739 ;
        RECT 60.464 19.278 60.51 36.248 ;
        RECT 43.536 36.206 60.464 36.294 ;
        RECT 48.136 31.606 65.065 31.693 ;
        RECT 60.418 19.324 60.464 36.294 ;
        RECT 43.49 36.252 60.418 36.34 ;
        RECT 48.182 31.56 65.111 31.647 ;
        RECT 60.372 19.37 60.418 36.34 ;
        RECT 43.444 36.298 60.372 36.386 ;
        RECT 48.228 31.514 65.157 31.601 ;
        RECT 60.326 19.416 60.372 36.386 ;
        RECT 43.398 36.344 60.326 36.432 ;
        RECT 48.274 31.468 65.203 31.555 ;
        RECT 60.28 19.462 60.326 36.432 ;
        RECT 43.352 36.39 60.28 36.478 ;
        RECT 48.32 31.422 65.249 31.509 ;
        RECT 60.234 19.508 60.28 36.478 ;
        RECT 43.306 36.436 60.234 36.524 ;
        RECT 48.366 31.376 65.295 31.463 ;
        RECT 60.188 19.554 60.234 36.524 ;
        RECT 43.26 36.482 60.188 36.57 ;
        RECT 48.412 31.33 65.341 31.417 ;
        RECT 60.142 19.6 60.188 36.57 ;
        RECT 43.214 36.528 60.142 36.616 ;
        RECT 48.458 31.284 65.387 31.371 ;
        RECT 60.096 19.646 60.142 36.616 ;
        RECT 43.168 36.574 60.096 36.662 ;
        RECT 48.504 31.238 65.433 31.325 ;
        RECT 60.05 19.692 60.096 36.662 ;
        RECT 43.122 36.62 60.05 36.708 ;
        RECT 48.55 31.192 65.479 31.279 ;
        RECT 60.004 19.738 60.05 36.708 ;
        RECT 43.076 36.666 60.004 36.754 ;
        RECT 48.596 31.146 65.525 31.233 ;
        RECT 59.958 19.784 60.004 36.754 ;
        RECT 43.03 36.712 59.958 36.8 ;
        RECT 48.642 31.1 65.571 31.187 ;
        RECT 59.912 19.83 59.958 36.8 ;
        RECT 42.984 36.758 59.912 36.846 ;
        RECT 48.688 31.054 65.617 31.141 ;
        RECT 59.866 19.876 59.912 36.846 ;
        RECT 42.938 36.804 59.866 36.892 ;
        RECT 48.734 31.008 65.663 31.095 ;
        RECT 59.82 19.922 59.866 36.892 ;
        RECT 42.892 36.85 59.82 36.938 ;
        RECT 48.78 30.962 65.709 31.049 ;
        RECT 59.774 19.968 59.82 36.938 ;
        RECT 42.846 36.896 59.774 36.984 ;
        RECT 48.826 30.916 65.755 31.003 ;
        RECT 59.728 20.014 59.774 36.984 ;
        RECT 42.8 36.942 59.728 37.03 ;
        RECT 48.872 30.87 65.801 30.957 ;
        RECT 59.682 20.06 59.728 37.03 ;
        RECT 42.754 36.988 59.682 37.076 ;
        RECT 48.918 30.824 65.847 30.911 ;
        RECT 59.636 20.106 59.682 37.076 ;
        RECT 42.708 37.034 59.636 37.122 ;
        RECT 48.964 30.778 65.893 30.865 ;
        RECT 59.59 20.152 59.636 37.122 ;
        RECT 42.662 37.08 59.59 37.168 ;
        RECT 49.01 30.732 65.939 30.819 ;
        RECT 59.544 20.198 59.59 37.168 ;
        RECT 42.616 37.126 59.544 37.214 ;
        RECT 49.056 30.686 65.985 30.773 ;
        RECT 59.498 20.244 59.544 37.214 ;
        RECT 42.57 37.172 59.498 37.26 ;
        RECT 49.102 30.64 66.031 30.727 ;
        RECT 59.452 20.29 59.498 37.26 ;
        RECT 42.524 37.218 59.452 37.306 ;
        RECT 49.148 30.594 66.077 30.681 ;
        RECT 59.406 20.336 59.452 37.306 ;
        RECT 42.478 37.264 59.406 37.352 ;
        RECT 49.194 30.548 66.123 30.635 ;
        RECT 59.36 20.382 59.406 37.352 ;
        RECT 42.432 37.31 59.36 37.398 ;
        RECT 49.24 30.502 66.169 30.589 ;
        RECT 59.314 20.428 59.36 37.398 ;
        RECT 42.386 37.356 59.314 37.444 ;
        RECT 49.286 30.456 66.215 30.543 ;
        RECT 59.268 20.474 59.314 37.444 ;
        RECT 42.34 37.402 59.268 37.49 ;
        RECT 49.332 30.41 66.261 30.497 ;
        RECT 59.222 20.52 59.268 37.49 ;
        RECT 42.294 37.448 59.222 37.536 ;
        RECT 49.378 30.364 66.307 30.451 ;
        RECT 59.176 20.566 59.222 37.536 ;
        RECT 42.248 37.494 59.176 37.582 ;
        RECT 49.424 30.318 66.353 30.405 ;
        RECT 59.13 20.612 59.176 37.582 ;
        RECT 42.202 37.54 59.13 37.628 ;
        RECT 49.47 30.272 66.399 30.359 ;
        RECT 59.084 20.658 59.13 37.628 ;
        RECT 42.156 37.586 59.084 37.674 ;
        RECT 49.516 30.226 66.445 30.313 ;
        RECT 59.038 20.704 59.084 37.674 ;
        RECT 42.11 37.632 59.038 37.72 ;
        RECT 49.562 30.18 66.491 30.267 ;
        RECT 58.992 20.75 59.038 37.72 ;
        RECT 42.064 37.678 58.992 37.766 ;
        RECT 49.608 30.134 66.537 30.221 ;
        RECT 58.946 20.796 58.992 37.766 ;
        RECT 42.018 37.724 58.946 37.812 ;
        RECT 49.654 30.088 66.583 30.175 ;
        RECT 58.9 20.842 58.946 37.812 ;
        RECT 41.972 37.77 58.9 37.858 ;
        RECT 49.7 30.042 66.629 30.129 ;
        RECT 58.854 20.888 58.9 37.858 ;
        RECT 41.926 37.816 58.854 37.904 ;
        RECT 49.746 29.996 66.675 30.083 ;
        RECT 58.808 20.934 58.854 37.904 ;
        RECT 41.88 37.862 58.808 37.95 ;
        RECT 49.792 29.95 66.721 30.037 ;
        RECT 58.762 20.98 58.808 37.95 ;
        RECT 41.834 37.908 58.762 37.996 ;
        RECT 49.838 29.904 66.767 29.991 ;
        RECT 58.716 21.026 58.762 37.996 ;
        RECT 41.788 37.954 58.716 38.042 ;
        RECT 49.884 29.858 66.813 29.945 ;
        RECT 58.67 21.072 58.716 38.042 ;
        RECT 41.742 38 58.67 38.088 ;
        RECT 49.93 29.812 66.859 29.899 ;
        RECT 58.624 21.118 58.67 38.088 ;
        RECT 41.696 38.046 58.624 38.134 ;
        RECT 49.976 29.766 66.905 29.853 ;
        RECT 58.578 21.164 58.624 38.134 ;
        RECT 41.65 38.092 58.578 38.18 ;
        RECT 50.022 29.72 66.951 29.807 ;
        RECT 58.532 21.21 58.578 38.18 ;
        RECT 41.604 38.138 58.532 38.226 ;
        RECT 50.068 29.674 66.997 29.761 ;
        RECT 58.486 21.256 58.532 38.226 ;
        RECT 41.558 38.184 58.486 38.272 ;
        RECT 50.114 29.628 67.043 29.715 ;
        RECT 58.44 21.302 58.486 38.272 ;
        RECT 41.512 38.23 58.44 38.318 ;
        RECT 50.16 29.582 67.089 29.669 ;
        RECT 58.394 21.348 58.44 38.318 ;
        RECT 41.466 38.276 58.394 38.364 ;
        RECT 50.206 29.536 67.135 29.623 ;
        RECT 58.348 21.394 58.394 38.364 ;
        RECT 41.42 38.322 58.348 38.41 ;
        RECT 50.252 29.49 67.181 29.577 ;
        RECT 58.302 21.44 58.348 38.41 ;
        RECT 41.374 38.368 58.302 38.456 ;
        RECT 50.298 29.444 67.227 29.531 ;
        RECT 58.256 21.486 58.302 38.456 ;
        RECT 41.328 38.414 58.256 38.502 ;
        RECT 50.344 29.398 67.273 29.485 ;
        RECT 58.21 21.532 58.256 38.502 ;
        RECT 41.282 38.46 58.21 38.548 ;
        RECT 50.39 29.352 67.319 29.439 ;
        RECT 58.164 21.578 58.21 38.548 ;
        RECT 41.236 38.506 58.164 38.594 ;
        RECT 50.436 29.306 67.365 29.393 ;
        RECT 58.118 21.624 58.164 38.594 ;
        RECT 41.19 38.552 58.118 38.64 ;
        RECT 50.482 29.26 67.411 29.347 ;
        RECT 58.072 21.67 58.118 38.64 ;
        RECT 41.144 38.598 58.072 38.686 ;
        RECT 50.528 29.214 67.457 29.301 ;
        RECT 58.026 21.716 58.072 38.686 ;
        RECT 41.098 38.644 58.026 38.732 ;
        RECT 50.574 29.168 67.503 29.255 ;
        RECT 57.98 21.762 58.026 38.732 ;
        RECT 41.052 38.69 57.98 38.778 ;
        RECT 50.62 29.122 67.549 29.209 ;
        RECT 57.934 21.808 57.98 38.778 ;
        RECT 41.006 38.736 57.934 38.824 ;
        RECT 50.666 29.076 67.595 29.163 ;
        RECT 57.888 21.854 57.934 38.824 ;
        RECT 40.96 38.782 57.888 38.87 ;
        RECT 50.712 29.03 67.641 29.117 ;
        RECT 57.842 21.9 57.888 38.87 ;
        RECT 40.914 38.828 57.842 38.916 ;
        RECT 50.758 28.984 67.687 29.071 ;
        RECT 57.796 21.946 57.842 38.916 ;
        RECT 40.868 38.874 57.796 38.962 ;
        RECT 50.804 28.938 110 29 ;
        RECT 57.75 21.992 57.796 38.962 ;
        RECT 40.822 38.92 57.75 39.008 ;
        RECT 50.85 28.892 110 29 ;
        RECT 57.704 22.038 57.75 39.008 ;
        RECT 40.776 38.966 57.704 39.054 ;
        RECT 50.896 28.846 110 29 ;
        RECT 57.658 22.084 57.704 39.054 ;
        RECT 40.73 39.012 57.658 39.1 ;
        RECT 50.942 28.8 110 29 ;
        RECT 57.612 22.13 57.658 39.1 ;
        RECT 40.684 39.058 57.612 39.146 ;
        RECT 50.988 28.754 110 29 ;
        RECT 57.566 22.176 57.612 39.146 ;
        RECT 40.638 39.104 57.566 39.192 ;
        RECT 51.034 28.708 110 29 ;
        RECT 57.52 22.222 57.566 39.192 ;
        RECT 40.592 39.15 57.52 39.238 ;
        RECT 51.08 28.662 110 29 ;
        RECT 57.474 22.268 57.52 39.238 ;
        RECT 40.546 39.196 57.474 39.284 ;
        RECT 51.126 28.616 110 29 ;
        RECT 57.428 22.314 57.474 39.284 ;
        RECT 40.5 39.242 57.428 39.33 ;
        RECT 51.172 28.57 110 29 ;
        RECT 57.382 22.36 57.428 39.33 ;
        RECT 40.454 39.288 57.382 39.376 ;
        RECT 51.218 28.524 110 29 ;
        RECT 57.336 22.406 57.382 39.376 ;
        RECT 40.408 39.334 57.336 39.422 ;
        RECT 51.264 28.478 110 29 ;
        RECT 57.29 22.452 57.336 39.422 ;
        RECT 40.362 39.38 57.29 39.468 ;
        RECT 51.31 28.432 110 29 ;
        RECT 57.244 22.498 57.29 39.468 ;
        RECT 40.316 39.426 57.244 39.514 ;
        RECT 51.356 28.386 110 29 ;
        RECT 57.198 22.544 57.244 39.514 ;
        RECT 40.27 39.472 57.198 39.56 ;
        RECT 51.402 28.34 110 29 ;
        RECT 57.152 22.59 57.198 39.56 ;
        RECT 40.224 39.518 57.152 39.606 ;
        RECT 51.448 28.294 110 29 ;
        RECT 57.106 22.636 57.152 39.606 ;
        RECT 40.178 39.564 57.106 39.652 ;
        RECT 51.494 28.248 110 29 ;
        RECT 57.06 22.682 57.106 39.652 ;
        RECT 40.132 39.61 57.06 39.698 ;
        RECT 51.54 28.202 110 29 ;
        RECT 57.014 22.728 57.06 39.698 ;
        RECT 40.086 39.656 57.014 39.744 ;
        RECT 51.586 28.156 110 29 ;
        RECT 56.968 22.774 57.014 39.744 ;
        RECT 40.04 39.702 56.968 39.79 ;
        RECT 51.632 28.11 110 29 ;
        RECT 56.922 22.82 56.968 39.79 ;
        RECT 39.994 39.748 56.922 39.836 ;
        RECT 51.678 28.064 110 29 ;
        RECT 56.876 22.866 56.922 39.836 ;
        RECT 39.948 39.794 56.876 39.882 ;
        RECT 51.724 28.018 110 29 ;
        RECT 56.83 22.912 56.876 39.882 ;
        RECT 39.902 39.84 56.83 39.928 ;
        RECT 51.77 27.972 110 29 ;
        RECT 56.784 22.958 56.83 39.928 ;
        RECT 39.856 39.886 56.784 39.974 ;
        RECT 51.816 27.926 110 29 ;
        RECT 56.738 23.004 56.784 39.974 ;
        RECT 39.81 39.932 56.738 40.02 ;
        RECT 51.862 27.88 110 29 ;
        RECT 56.692 23.05 56.738 40.02 ;
        RECT 39.764 39.978 56.692 40.066 ;
        RECT 51.908 27.834 110 29 ;
        RECT 56.646 23.096 56.692 40.066 ;
        RECT 39.718 40.024 56.646 40.112 ;
        RECT 51.954 27.788 110 29 ;
        RECT 56.6 23.142 56.646 40.112 ;
        RECT 39.672 40.07 56.6 40.158 ;
        RECT 52 27.742 110 29 ;
        RECT 56.554 23.188 56.6 40.158 ;
        RECT 39.626 40.116 56.554 40.204 ;
        RECT 52.046 27.696 110 29 ;
        RECT 56.508 23.234 56.554 40.204 ;
        RECT 39.58 40.162 56.508 40.25 ;
        RECT 52.092 27.65 110 29 ;
        RECT 56.462 23.28 56.508 40.25 ;
        RECT 39.534 40.208 56.462 40.296 ;
        RECT 52.138 27.604 110 29 ;
        RECT 56.416 23.326 56.462 40.296 ;
        RECT 39.488 40.254 56.416 40.342 ;
        RECT 52.184 27.558 110 29 ;
        RECT 56.37 23.372 56.416 40.342 ;
        RECT 39.442 40.3 56.37 40.388 ;
        RECT 52.23 27.512 110 29 ;
        RECT 56.324 23.418 56.37 40.388 ;
        RECT 39.396 40.346 56.324 40.434 ;
        RECT 52.276 27.466 110 29 ;
        RECT 56.278 23.464 56.324 40.434 ;
        RECT 39.35 40.392 56.278 40.48 ;
        RECT 52.322 27.42 110 29 ;
        RECT 56.232 23.51 56.278 40.48 ;
        RECT 39.304 40.438 56.232 40.526 ;
        RECT 52.368 27.374 110 29 ;
        RECT 56.186 23.556 56.232 40.526 ;
        RECT 39.258 40.484 56.186 40.572 ;
        RECT 52.414 27.328 110 29 ;
        RECT 56.14 23.602 56.186 40.572 ;
        RECT 39.212 40.53 56.14 40.618 ;
        RECT 52.46 27.282 110 29 ;
        RECT 56.094 23.648 56.14 40.618 ;
        RECT 39.166 40.576 56.094 40.664 ;
        RECT 52.506 27.236 110 29 ;
        RECT 56.048 23.694 56.094 40.664 ;
        RECT 39.12 40.622 56.048 40.71 ;
        RECT 52.552 27.19 110 29 ;
        RECT 56.002 23.74 56.048 40.71 ;
        RECT 39.074 40.668 56.002 40.756 ;
        RECT 52.598 27.144 110 29 ;
        RECT 55.956 23.786 56.002 40.756 ;
        RECT 39.028 40.714 55.956 40.802 ;
        RECT 52.644 27.098 110 29 ;
        RECT 55.91 23.832 55.956 40.802 ;
        RECT 38.982 40.76 55.91 40.848 ;
        RECT 52.69 27.052 110 29 ;
        RECT 55.864 23.878 55.91 40.848 ;
        RECT 38.936 40.806 55.864 40.894 ;
        RECT 52.736 27.006 110 29 ;
        RECT 55.818 23.924 55.864 40.894 ;
        RECT 38.89 40.852 55.818 40.94 ;
        RECT 52.782 26.96 110 29 ;
        RECT 55.772 23.97 55.818 40.94 ;
        RECT 38.844 40.898 55.772 40.986 ;
        RECT 52.828 26.914 110 29 ;
        RECT 55.726 24.016 55.772 40.986 ;
        RECT 38.798 40.944 55.726 41.032 ;
        RECT 52.874 26.868 110 29 ;
        RECT 55.68 24.062 55.726 41.032 ;
        RECT 38.752 40.99 55.68 41.078 ;
        RECT 52.92 26.822 110 29 ;
        RECT 55.634 24.108 55.68 41.078 ;
        RECT 38.706 41.036 55.634 41.124 ;
        RECT 52.966 26.776 110 29 ;
        RECT 55.588 24.154 55.634 41.124 ;
        RECT 38.66 41.082 55.588 41.17 ;
        RECT 53.012 26.73 110 29 ;
        RECT 55.542 24.2 55.588 41.17 ;
        RECT 38.614 41.128 55.542 41.216 ;
        RECT 53.058 26.684 110 29 ;
        RECT 55.496 24.246 55.542 41.216 ;
        RECT 38.568 41.174 55.496 41.262 ;
        RECT 53.104 26.638 110 29 ;
        RECT 55.45 24.292 55.496 41.262 ;
        RECT 38.522 41.22 55.45 41.308 ;
        RECT 53.15 26.592 110 29 ;
        RECT 55.404 24.338 55.45 41.308 ;
        RECT 38.476 41.266 55.404 41.354 ;
        RECT 53.196 26.546 110 29 ;
        RECT 55.358 24.384 55.404 41.354 ;
        RECT 38.43 41.312 55.358 41.4 ;
        RECT 53.242 26.5 110 29 ;
        RECT 55.312 24.43 55.358 41.4 ;
        RECT 38.384 41.358 55.312 41.446 ;
        RECT 53.288 26.454 110 29 ;
        RECT 55.266 24.476 55.312 41.446 ;
        RECT 38.338 41.404 55.266 41.492 ;
        RECT 53.334 26.408 110 29 ;
        RECT 55.22 24.522 55.266 41.492 ;
        RECT 38.292 41.45 55.22 41.538 ;
        RECT 53.38 26.362 110 29 ;
        RECT 55.174 24.568 55.22 41.538 ;
        RECT 38.246 41.496 55.174 41.584 ;
        RECT 53.426 26.316 110 29 ;
        RECT 55.128 24.614 55.174 41.584 ;
        RECT 38.2 41.542 55.128 41.63 ;
        RECT 53.472 26.27 110 29 ;
        RECT 55.082 24.66 55.128 41.63 ;
        RECT 38.154 41.588 55.082 41.676 ;
        RECT 53.518 26.224 110 29 ;
        RECT 55.036 24.706 55.082 41.676 ;
        RECT 38.108 41.634 55.036 41.722 ;
        RECT 53.564 26.178 110 29 ;
        RECT 54.99 24.752 55.036 41.722 ;
        RECT 38.062 41.68 54.99 41.768 ;
        RECT 53.61 26.132 110 29 ;
        RECT 54.944 24.798 54.99 41.768 ;
        RECT 38.016 41.726 54.944 41.814 ;
        RECT 53.656 26.086 110 29 ;
        RECT 54.898 24.844 54.944 41.814 ;
        RECT 37.97 41.772 54.898 41.86 ;
        RECT 53.702 26.04 110 29 ;
        RECT 54.852 24.89 54.898 41.86 ;
        RECT 37.924 41.818 54.852 41.906 ;
        RECT 53.748 25.994 110 29 ;
        RECT 54.806 24.936 54.852 41.906 ;
        RECT 37.878 41.864 54.806 41.952 ;
        RECT 53.794 25.948 110 29 ;
        RECT 54.76 24.982 54.806 41.952 ;
        RECT 37.832 41.91 54.76 41.998 ;
        RECT 53.84 25.902 110 29 ;
        RECT 54.714 25.028 54.76 41.998 ;
        RECT 37.786 41.956 54.714 42.044 ;
        RECT 53.886 25.856 110 29 ;
        RECT 54.668 25.074 54.714 42.044 ;
        RECT 37.74 42.002 54.668 42.09 ;
        RECT 53.932 25.81 110 29 ;
        RECT 54.622 25.12 54.668 42.09 ;
        RECT 37.694 42.048 54.622 42.136 ;
        RECT 53.978 25.764 110 29 ;
        RECT 54.576 25.166 54.622 42.136 ;
        RECT 37.648 42.094 54.576 42.182 ;
        RECT 54.024 25.718 110 29 ;
        RECT 54.53 25.212 54.576 42.182 ;
        RECT 37.602 42.14 54.53 42.228 ;
        RECT 54.07 25.672 110 29 ;
        RECT 54.484 25.258 54.53 42.228 ;
        RECT 37.556 42.186 54.484 42.274 ;
        RECT 54.116 25.626 110 29 ;
        RECT 54.438 25.304 54.484 42.274 ;
        RECT 37.51 42.232 54.438 42.32 ;
        RECT 54.162 25.58 110 29 ;
        RECT 54.392 25.35 54.438 42.32 ;
        RECT 37.464 42.278 54.392 42.366 ;
        RECT 54.208 25.534 110 29 ;
        RECT 54.346 25.396 54.392 42.366 ;
        RECT 37.418 42.324 54.346 42.412 ;
        RECT 54.254 25.488 110 29 ;
        RECT 54.3 25.442 54.346 42.412 ;
        RECT 37.372 42.37 54.3 42.458 ;
        RECT 37.326 42.416 54.254 42.504 ;
        RECT 37.28 42.462 54.208 42.55 ;
        RECT 37.234 42.508 54.162 42.596 ;
        RECT 37.188 42.554 54.116 42.642 ;
        RECT 37.142 42.6 54.07 42.688 ;
        RECT 37.096 42.646 54.024 42.734 ;
        RECT 37.05 42.692 53.978 42.78 ;
        RECT 37.004 42.738 53.932 42.826 ;
        RECT 36.958 42.784 53.886 42.872 ;
        RECT 36.912 42.83 53.84 42.918 ;
        RECT 36.866 42.876 53.794 42.964 ;
        RECT 36.82 42.922 53.748 43.01 ;
        RECT 36.774 42.968 53.702 43.056 ;
        RECT 36.728 43.014 53.656 43.102 ;
        RECT 36.682 43.06 53.61 43.148 ;
        RECT 36.636 43.106 53.564 43.194 ;
        RECT 36.59 43.152 53.518 43.24 ;
        RECT 36.544 43.198 53.472 43.286 ;
        RECT 36.498 43.244 53.426 43.332 ;
        RECT 36.452 43.29 53.38 43.378 ;
        RECT 36.406 43.336 53.334 43.424 ;
        RECT 36.36 43.382 53.288 43.47 ;
        RECT 36.314 43.428 53.242 43.516 ;
        RECT 36.268 43.474 53.196 43.562 ;
        RECT 36.222 43.52 53.15 43.608 ;
        RECT 36.176 43.566 53.104 43.654 ;
        RECT 36.13 43.612 53.058 43.7 ;
        RECT 36.084 43.658 53.012 43.746 ;
        RECT 36.038 43.704 52.966 43.792 ;
        RECT 35.992 43.75 52.92 43.838 ;
        RECT 35.946 43.796 52.874 43.884 ;
        RECT 35.9 43.842 52.828 43.93 ;
        RECT 35.854 43.888 52.782 43.976 ;
        RECT 35.808 43.934 52.736 44.022 ;
        RECT 35.762 43.98 52.69 44.068 ;
        RECT 35.716 44.026 52.644 44.114 ;
        RECT 35.67 44.072 52.598 44.16 ;
        RECT 35.624 44.118 52.552 44.206 ;
        RECT 35.578 44.164 52.506 44.252 ;
        RECT 35.532 44.21 52.46 44.298 ;
        RECT 35.486 44.256 52.414 44.344 ;
        RECT 35.44 44.302 52.368 44.39 ;
        RECT 35.394 44.348 52.322 44.436 ;
        RECT 35.348 44.394 52.276 44.482 ;
        RECT 35.302 44.44 52.23 44.528 ;
        RECT 35.256 44.486 52.184 44.574 ;
        RECT 35.21 44.532 52.138 44.62 ;
        RECT 35.164 44.578 52.092 44.666 ;
        RECT 35.118 44.624 52.046 44.712 ;
        RECT 35.072 44.67 52 44.758 ;
        RECT 35.026 44.716 51.954 44.804 ;
        RECT 34.98 44.762 51.908 44.85 ;
        RECT 34.934 44.808 51.862 44.896 ;
        RECT 34.888 44.854 51.816 44.942 ;
        RECT 34.842 44.9 51.77 44.988 ;
        RECT 34.796 44.946 51.724 45.034 ;
        RECT 34.75 44.992 51.678 45.08 ;
        RECT 34.704 45.038 51.632 45.126 ;
        RECT 34.658 45.084 51.586 45.172 ;
        RECT 34.612 45.13 51.54 45.218 ;
        RECT 34.566 45.176 51.494 45.264 ;
        RECT 34.52 45.222 51.448 45.31 ;
        RECT 34.474 45.268 51.402 45.356 ;
        RECT 34.428 45.314 51.356 45.402 ;
        RECT 34.382 45.36 51.31 45.448 ;
        RECT 34.336 45.406 51.264 45.494 ;
        RECT 34.29 45.452 51.218 45.54 ;
        RECT 34.244 45.498 51.172 45.586 ;
        RECT 34.198 45.544 51.126 45.632 ;
        RECT 34.152 45.59 51.08 45.678 ;
        RECT 34.106 45.636 51.034 45.724 ;
        RECT 34.06 45.682 50.988 45.77 ;
        RECT 34.014 45.728 50.942 45.816 ;
        RECT 33.968 45.774 50.896 45.862 ;
        RECT 33.922 45.82 50.85 45.908 ;
        RECT 33.876 45.866 50.804 45.954 ;
        RECT 33.83 45.912 50.758 46 ;
        RECT 33.784 45.958 50.712 46.046 ;
        RECT 33.738 46.004 50.666 46.092 ;
        RECT 33.692 46.05 50.62 46.138 ;
        RECT 33.646 46.096 50.574 46.184 ;
        RECT 33.6 46.142 50.528 46.23 ;
        RECT 33.554 46.188 50.482 46.276 ;
        RECT 33.508 46.234 50.436 46.322 ;
        RECT 33.462 46.28 50.39 46.368 ;
        RECT 33.416 46.326 50.344 46.414 ;
        RECT 33.37 46.372 50.298 46.46 ;
        RECT 33.324 46.418 50.252 46.506 ;
        RECT 33.278 46.464 50.206 46.552 ;
        RECT 33.232 46.51 50.16 46.598 ;
        RECT 33.186 46.556 50.114 46.644 ;
        RECT 33.14 46.602 50.068 46.69 ;
        RECT 33.094 46.648 50.022 46.736 ;
        RECT 33.048 46.694 49.976 46.782 ;
        RECT 33.002 46.74 49.93 46.828 ;
        RECT 32.956 46.786 49.884 46.874 ;
        RECT 32.91 46.832 49.838 46.92 ;
        RECT 32.864 46.878 49.792 46.966 ;
        RECT 32.818 46.924 49.746 47.012 ;
        RECT 32.772 46.97 49.7 47.058 ;
        RECT 32.726 47.016 49.654 47.104 ;
        RECT 32.68 47.062 49.608 47.15 ;
        RECT 32.634 47.108 49.562 47.196 ;
        RECT 32.588 47.154 49.516 47.242 ;
        RECT 32.542 47.2 49.47 47.288 ;
        RECT 32.496 47.246 49.424 47.334 ;
        RECT 32.45 47.292 49.378 47.38 ;
        RECT 32.404 47.338 49.332 47.426 ;
        RECT 32.358 47.384 49.286 47.472 ;
        RECT 32.312 47.43 49.24 47.518 ;
        RECT 32.266 47.476 49.194 47.564 ;
        RECT 32.22 47.522 49.148 47.61 ;
        RECT 32.174 47.568 49.102 47.656 ;
        RECT 32.128 47.614 49.056 47.702 ;
        RECT 32.082 47.66 49.01 47.748 ;
        RECT 32.036 47.706 48.964 47.794 ;
        RECT 31.99 47.752 48.918 47.84 ;
        RECT 31.944 47.798 48.872 47.886 ;
        RECT 31.898 47.844 48.826 47.932 ;
        RECT 31.852 47.89 48.78 47.978 ;
        RECT 31.806 47.936 48.734 48.024 ;
        RECT 31.76 47.982 48.688 48.07 ;
        RECT 31.714 48.028 48.642 48.116 ;
        RECT 31.668 48.074 48.596 48.162 ;
        RECT 31.622 48.12 48.55 48.208 ;
        RECT 31.576 48.166 48.504 48.254 ;
        RECT 31.53 48.212 48.458 48.3 ;
        RECT 31.484 48.258 48.412 48.346 ;
        RECT 31.438 48.304 48.366 48.392 ;
        RECT 31.392 48.35 48.32 48.438 ;
        RECT 31.346 48.396 48.274 48.484 ;
        RECT 31.3 48.442 48.228 48.53 ;
        RECT 31.254 48.488 48.182 48.576 ;
        RECT 31.208 48.534 48.136 48.622 ;
        RECT 31.162 48.58 48.09 48.668 ;
        RECT 31.116 48.626 48.044 48.714 ;
        RECT 31.07 48.672 47.998 48.76 ;
        RECT 31.024 48.718 47.952 48.806 ;
        RECT 30.978 48.764 47.906 48.852 ;
        RECT 30.932 48.81 47.86 48.898 ;
        RECT 30.886 48.856 47.814 48.944 ;
        RECT 30.84 48.902 47.768 48.99 ;
        RECT 30.794 48.948 47.722 49.036 ;
        RECT 30.748 48.994 47.676 49.082 ;
        RECT 30.702 49.04 47.63 49.128 ;
        RECT 30.656 49.086 47.584 49.174 ;
        RECT 30.61 49.132 47.538 49.22 ;
        RECT 30.564 49.178 47.492 49.266 ;
        RECT 30.518 49.224 47.446 49.312 ;
        RECT 30.472 49.27 47.4 49.358 ;
        RECT 30.426 49.316 47.354 49.404 ;
        RECT 30.38 49.362 47.308 49.45 ;
        RECT 30.334 49.408 47.262 49.496 ;
        RECT 30.288 49.454 47.216 49.542 ;
        RECT 30.242 49.5 47.17 49.588 ;
        RECT 30.196 49.546 47.124 49.634 ;
        RECT 30.15 49.592 47.078 49.68 ;
        RECT 30.104 49.638 47.032 49.726 ;
        RECT 30.058 49.684 46.986 49.772 ;
        RECT 30.012 49.73 46.94 49.818 ;
        RECT 29.966 49.776 46.894 49.864 ;
        RECT 29.92 49.822 46.848 49.91 ;
        RECT 29.874 49.868 46.802 49.956 ;
        RECT 29.828 49.914 46.756 50.002 ;
        RECT 29.782 49.96 46.71 50.048 ;
        RECT 29.736 50.006 46.664 50.094 ;
        RECT 29.69 50.052 46.618 50.14 ;
        RECT 29.644 50.098 46.572 50.186 ;
        RECT 29.598 50.144 46.526 50.232 ;
        RECT 29.552 50.19 46.48 50.278 ;
        RECT 29.506 50.236 46.434 50.324 ;
        RECT 29.46 50.282 46.388 50.37 ;
        RECT 29.414 50.328 46.342 50.416 ;
        RECT 29.368 50.374 46.296 50.462 ;
        RECT 29.322 50.42 46.25 50.508 ;
        RECT 29.276 50.466 46.204 50.554 ;
        RECT 29.23 50.512 46.158 50.6 ;
        RECT 29.184 50.558 46.112 50.646 ;
        RECT 29.138 50.604 46.066 50.692 ;
        RECT 29.092 50.65 46.02 50.738 ;
        RECT 29 50.742 45.974 50.784 ;
        RECT 29.046 50.696 45.974 50.784 ;
        RECT 28.96 50.785 45.928 50.83 ;
        RECT 28.914 50.828 45.882 50.876 ;
        RECT 28.868 50.874 45.836 50.922 ;
        RECT 28.822 50.92 45.79 50.968 ;
        RECT 28.776 50.966 45.744 51.014 ;
        RECT 28.73 51.012 45.698 51.06 ;
        RECT 28.684 51.058 45.652 51.106 ;
        RECT 28.638 51.104 45.606 51.152 ;
        RECT 28.592 51.15 45.56 51.198 ;
        RECT 28.546 51.196 45.514 51.244 ;
        RECT 28.5 51.242 45.468 51.29 ;
        RECT 28.454 51.288 45.422 51.336 ;
        RECT 28.408 51.334 45.376 51.382 ;
        RECT 56.015 3.5 110 15.5 ;
        RECT 39.052 20.44 56.015 20.488 ;
        RECT 39.098 20.394 56.061 20.447 ;
        RECT 55.98 3.517 56.015 20.488 ;
        RECT 39.144 20.348 56.107 20.401 ;
        RECT 55.934 3.558 55.98 20.528 ;
        RECT 39.006 20.486 55.934 20.574 ;
        RECT 39.19 20.302 56.153 20.355 ;
        RECT 55.888 3.604 55.934 20.574 ;
        RECT 38.96 20.532 55.888 20.62 ;
        RECT 39.236 20.256 56.199 20.309 ;
        RECT 55.842 3.65 55.888 20.62 ;
        RECT 38.914 20.578 55.842 20.666 ;
        RECT 39.282 20.21 56.245 20.263 ;
        RECT 55.796 3.696 55.842 20.666 ;
        RECT 38.868 20.624 55.796 20.712 ;
        RECT 39.328 20.164 56.291 20.217 ;
        RECT 55.75 3.742 55.796 20.712 ;
        RECT 38.822 20.67 55.75 20.758 ;
        RECT 39.374 20.118 56.337 20.171 ;
        RECT 55.704 3.788 55.75 20.758 ;
        RECT 38.776 20.716 55.704 20.804 ;
        RECT 39.42 20.072 56.383 20.125 ;
        RECT 55.658 3.834 55.704 20.804 ;
        RECT 38.73 20.762 55.658 20.85 ;
        RECT 39.466 20.026 56.429 20.079 ;
        RECT 55.612 3.88 55.658 20.85 ;
        RECT 38.684 20.808 55.612 20.896 ;
        RECT 39.512 19.98 56.475 20.033 ;
        RECT 55.566 3.926 55.612 20.896 ;
        RECT 38.638 20.854 55.566 20.942 ;
        RECT 39.558 19.934 56.521 19.987 ;
        RECT 55.52 3.972 55.566 20.942 ;
        RECT 38.592 20.9 55.52 20.988 ;
        RECT 39.604 19.888 56.567 19.941 ;
        RECT 55.474 4.018 55.52 20.988 ;
        RECT 38.546 20.946 55.474 21.034 ;
        RECT 39.65 19.842 56.613 19.895 ;
        RECT 55.428 4.064 55.474 21.034 ;
        RECT 38.5 20.992 55.428 21.08 ;
        RECT 39.696 19.796 56.659 19.849 ;
        RECT 55.382 4.11 55.428 21.08 ;
        RECT 38.454 21.038 55.382 21.126 ;
        RECT 39.742 19.75 56.705 19.803 ;
        RECT 55.336 4.156 55.382 21.126 ;
        RECT 38.408 21.084 55.336 21.172 ;
        RECT 39.788 19.704 56.751 19.757 ;
        RECT 55.29 4.202 55.336 21.172 ;
        RECT 38.362 21.13 55.29 21.218 ;
        RECT 39.834 19.658 56.797 19.711 ;
        RECT 55.244 4.248 55.29 21.218 ;
        RECT 38.316 21.176 55.244 21.264 ;
        RECT 39.88 19.612 56.843 19.665 ;
        RECT 55.198 4.294 55.244 21.264 ;
        RECT 38.27 21.222 55.198 21.31 ;
        RECT 39.926 19.566 56.889 19.619 ;
        RECT 55.152 4.34 55.198 21.31 ;
        RECT 38.224 21.268 55.152 21.356 ;
        RECT 39.972 19.52 56.935 19.573 ;
        RECT 55.106 4.386 55.152 21.356 ;
        RECT 38.178 21.314 55.106 21.402 ;
        RECT 40.018 19.474 56.981 19.527 ;
        RECT 55.06 4.432 55.106 21.402 ;
        RECT 38.132 21.36 55.06 21.448 ;
        RECT 40.064 19.428 57.027 19.481 ;
        RECT 55.014 4.478 55.06 21.448 ;
        RECT 38.086 21.406 55.014 21.494 ;
        RECT 40.11 19.382 57.073 19.435 ;
        RECT 54.968 4.524 55.014 21.494 ;
        RECT 38.04 21.452 54.968 21.54 ;
        RECT 40.156 19.336 57.119 19.389 ;
        RECT 54.922 4.57 54.968 21.54 ;
        RECT 37.994 21.498 54.922 21.586 ;
        RECT 40.202 19.29 57.165 19.343 ;
        RECT 54.876 4.616 54.922 21.586 ;
        RECT 37.948 21.544 54.876 21.632 ;
        RECT 40.248 19.244 57.211 19.297 ;
        RECT 54.83 4.662 54.876 21.632 ;
        RECT 37.902 21.59 54.83 21.678 ;
        RECT 40.294 19.198 57.257 19.251 ;
        RECT 54.784 4.708 54.83 21.678 ;
        RECT 37.856 21.636 54.784 21.724 ;
        RECT 40.34 19.152 57.303 19.205 ;
        RECT 54.738 4.754 54.784 21.724 ;
        RECT 37.81 21.682 54.738 21.77 ;
        RECT 40.386 19.106 57.349 19.159 ;
        RECT 54.692 4.8 54.738 21.77 ;
        RECT 37.764 21.728 54.692 21.816 ;
        RECT 40.432 19.06 57.395 19.113 ;
        RECT 54.646 4.846 54.692 21.816 ;
        RECT 37.718 21.774 54.646 21.862 ;
        RECT 40.478 19.014 57.441 19.067 ;
        RECT 54.6 4.892 54.646 21.862 ;
        RECT 37.672 21.82 54.6 21.908 ;
        RECT 40.524 18.968 57.487 19.021 ;
        RECT 54.554 4.938 54.6 21.908 ;
        RECT 37.626 21.866 54.554 21.954 ;
        RECT 40.57 18.922 57.533 18.975 ;
        RECT 54.508 4.984 54.554 21.954 ;
        RECT 37.58 21.912 54.508 22 ;
        RECT 40.616 18.876 57.579 18.929 ;
        RECT 54.462 5.03 54.508 22 ;
        RECT 37.534 21.958 54.462 22.046 ;
        RECT 40.662 18.83 57.625 18.883 ;
        RECT 54.416 5.076 54.462 22.046 ;
        RECT 37.488 22.004 54.416 22.092 ;
        RECT 40.708 18.784 57.671 18.837 ;
        RECT 54.37 5.122 54.416 22.092 ;
        RECT 37.442 22.05 54.37 22.138 ;
        RECT 40.754 18.738 57.717 18.791 ;
        RECT 54.324 5.168 54.37 22.138 ;
        RECT 37.396 22.096 54.324 22.184 ;
        RECT 40.8 18.692 57.763 18.745 ;
        RECT 54.278 5.214 54.324 22.184 ;
        RECT 37.35 22.142 54.278 22.23 ;
        RECT 40.846 18.646 57.809 18.699 ;
        RECT 54.232 5.26 54.278 22.23 ;
        RECT 37.304 22.188 54.232 22.276 ;
        RECT 40.892 18.6 57.855 18.653 ;
        RECT 54.186 5.306 54.232 22.276 ;
        RECT 37.258 22.234 54.186 22.322 ;
        RECT 40.938 18.554 57.901 18.607 ;
        RECT 54.14 5.352 54.186 22.322 ;
        RECT 37.212 22.28 54.14 22.368 ;
        RECT 40.984 18.508 57.947 18.561 ;
        RECT 54.094 5.398 54.14 22.368 ;
        RECT 37.166 22.326 54.094 22.414 ;
        RECT 41.03 18.462 57.993 18.515 ;
        RECT 54.048 5.444 54.094 22.414 ;
        RECT 37.12 22.372 54.048 22.46 ;
        RECT 41.076 18.416 58.039 18.469 ;
        RECT 54.002 5.49 54.048 22.46 ;
        RECT 37.074 22.418 54.002 22.506 ;
        RECT 41.122 18.37 58.085 18.423 ;
        RECT 53.956 5.536 54.002 22.506 ;
        RECT 37.028 22.464 53.956 22.552 ;
        RECT 41.168 18.324 58.131 18.377 ;
        RECT 53.91 5.582 53.956 22.552 ;
        RECT 36.982 22.51 53.91 22.598 ;
        RECT 41.214 18.278 58.177 18.331 ;
        RECT 53.864 5.628 53.91 22.598 ;
        RECT 36.936 22.556 53.864 22.644 ;
        RECT 41.26 18.232 58.223 18.285 ;
        RECT 53.818 5.674 53.864 22.644 ;
        RECT 36.89 22.602 53.818 22.69 ;
        RECT 41.306 18.186 58.269 18.239 ;
        RECT 53.772 5.72 53.818 22.69 ;
        RECT 36.844 22.648 53.772 22.736 ;
        RECT 41.352 18.14 58.315 18.193 ;
        RECT 53.726 5.766 53.772 22.736 ;
        RECT 36.798 22.694 53.726 22.782 ;
        RECT 41.398 18.094 58.361 18.147 ;
        RECT 53.68 5.812 53.726 22.782 ;
        RECT 36.752 22.74 53.68 22.828 ;
        RECT 41.444 18.048 58.407 18.101 ;
        RECT 53.634 5.858 53.68 22.828 ;
        RECT 36.706 22.786 53.634 22.874 ;
        RECT 41.49 18.002 58.453 18.055 ;
        RECT 53.588 5.904 53.634 22.874 ;
        RECT 36.66 22.832 53.588 22.92 ;
        RECT 41.536 17.956 58.499 18.009 ;
        RECT 53.542 5.95 53.588 22.92 ;
        RECT 36.614 22.878 53.542 22.966 ;
        RECT 41.582 17.91 58.545 17.963 ;
        RECT 53.496 5.996 53.542 22.966 ;
        RECT 36.568 22.924 53.496 23.012 ;
        RECT 41.628 17.864 58.591 17.917 ;
        RECT 53.45 6.042 53.496 23.012 ;
        RECT 36.522 22.97 53.45 23.058 ;
        RECT 41.674 17.818 58.637 17.871 ;
        RECT 53.404 6.088 53.45 23.058 ;
        RECT 36.476 23.016 53.404 23.104 ;
        RECT 41.72 17.772 58.683 17.825 ;
        RECT 53.358 6.134 53.404 23.104 ;
        RECT 36.43 23.062 53.358 23.15 ;
        RECT 41.766 17.726 58.729 17.779 ;
        RECT 53.312 6.18 53.358 23.15 ;
        RECT 36.384 23.108 53.312 23.196 ;
        RECT 41.812 17.68 58.775 17.733 ;
        RECT 53.266 6.226 53.312 23.196 ;
        RECT 36.338 23.154 53.266 23.242 ;
        RECT 41.858 17.634 58.821 17.687 ;
        RECT 53.22 6.272 53.266 23.242 ;
        RECT 36.292 23.2 53.22 23.288 ;
        RECT 41.904 17.588 58.867 17.641 ;
        RECT 53.174 6.318 53.22 23.288 ;
        RECT 36.246 23.246 53.174 23.334 ;
        RECT 41.95 17.542 58.913 17.595 ;
        RECT 53.128 6.364 53.174 23.334 ;
        RECT 36.2 23.292 53.128 23.38 ;
        RECT 41.996 17.496 58.959 17.549 ;
        RECT 53.082 6.41 53.128 23.38 ;
        RECT 36.154 23.338 53.082 23.426 ;
        RECT 42.042 17.45 59.005 17.503 ;
        RECT 53.036 6.456 53.082 23.426 ;
        RECT 36.108 23.384 53.036 23.472 ;
        RECT 42.088 17.404 59.051 17.457 ;
        RECT 52.99 6.502 53.036 23.472 ;
        RECT 36.062 23.43 52.99 23.518 ;
        RECT 42.134 17.358 59.097 17.411 ;
        RECT 52.944 6.548 52.99 23.518 ;
        RECT 36.016 23.476 52.944 23.564 ;
        RECT 42.18 17.312 59.143 17.365 ;
        RECT 52.898 6.594 52.944 23.564 ;
        RECT 35.97 23.522 52.898 23.61 ;
        RECT 42.226 17.266 59.189 17.319 ;
        RECT 52.852 6.64 52.898 23.61 ;
        RECT 35.924 23.568 52.852 23.656 ;
        RECT 42.272 17.22 59.235 17.273 ;
        RECT 52.806 6.686 52.852 23.656 ;
        RECT 35.878 23.614 52.806 23.702 ;
        RECT 42.318 17.174 59.281 17.227 ;
        RECT 52.76 6.732 52.806 23.702 ;
        RECT 35.832 23.66 52.76 23.748 ;
        RECT 42.364 17.128 59.327 17.181 ;
        RECT 52.714 6.778 52.76 23.748 ;
        RECT 35.786 23.706 52.714 23.794 ;
        RECT 42.41 17.082 59.373 17.135 ;
        RECT 52.668 6.824 52.714 23.794 ;
        RECT 35.74 23.752 52.668 23.84 ;
        RECT 42.456 17.036 59.419 17.089 ;
        RECT 52.622 6.87 52.668 23.84 ;
        RECT 35.694 23.798 52.622 23.886 ;
        RECT 42.502 16.99 59.465 17.043 ;
        RECT 52.576 6.916 52.622 23.886 ;
        RECT 35.648 23.844 52.576 23.932 ;
        RECT 42.548 16.944 59.511 16.997 ;
        RECT 52.53 6.962 52.576 23.932 ;
        RECT 35.602 23.89 52.53 23.978 ;
        RECT 42.594 16.898 59.557 16.951 ;
        RECT 52.484 7.008 52.53 23.978 ;
        RECT 35.556 23.936 52.484 24.024 ;
        RECT 42.64 16.852 59.603 16.905 ;
        RECT 52.438 7.054 52.484 24.024 ;
        RECT 35.51 23.982 52.438 24.07 ;
        RECT 42.686 16.806 59.649 16.859 ;
        RECT 52.392 7.1 52.438 24.07 ;
        RECT 35.464 24.028 52.392 24.116 ;
        RECT 42.732 16.76 59.695 16.813 ;
        RECT 52.346 7.146 52.392 24.116 ;
        RECT 35.418 24.074 52.346 24.162 ;
        RECT 42.778 16.714 59.741 16.767 ;
        RECT 52.3 7.192 52.346 24.162 ;
        RECT 35.372 24.12 52.3 24.208 ;
        RECT 42.824 16.668 59.787 16.721 ;
        RECT 52.254 7.238 52.3 24.208 ;
        RECT 35.326 24.166 52.254 24.254 ;
        RECT 42.87 16.622 59.833 16.675 ;
        RECT 52.208 7.284 52.254 24.254 ;
        RECT 35.28 24.212 52.208 24.3 ;
        RECT 42.916 16.576 59.879 16.629 ;
        RECT 52.162 7.33 52.208 24.3 ;
        RECT 35.234 24.258 52.162 24.346 ;
        RECT 42.962 16.53 59.925 16.583 ;
        RECT 52.116 7.376 52.162 24.346 ;
        RECT 35.188 24.304 52.116 24.392 ;
        RECT 43.008 16.484 59.971 16.537 ;
        RECT 52.07 7.422 52.116 24.392 ;
        RECT 35.142 24.35 52.07 24.438 ;
        RECT 43.054 16.438 60.017 16.491 ;
        RECT 52.024 7.468 52.07 24.438 ;
        RECT 35.096 24.396 52.024 24.484 ;
        RECT 43.1 16.392 60.063 16.445 ;
        RECT 51.978 7.514 52.024 24.484 ;
        RECT 35.05 24.442 51.978 24.53 ;
        RECT 43.146 16.346 60.109 16.399 ;
        RECT 51.932 7.56 51.978 24.53 ;
        RECT 35.004 24.488 51.932 24.576 ;
        RECT 43.192 16.3 60.155 16.353 ;
        RECT 51.886 7.606 51.932 24.576 ;
        RECT 34.958 24.534 51.886 24.622 ;
        RECT 43.238 16.254 60.201 16.307 ;
        RECT 51.84 7.652 51.886 24.622 ;
        RECT 34.912 24.58 51.84 24.668 ;
        RECT 43.284 16.208 60.247 16.261 ;
        RECT 51.794 7.698 51.84 24.668 ;
        RECT 34.866 24.626 51.794 24.714 ;
        RECT 43.33 16.162 60.293 16.215 ;
        RECT 51.748 7.744 51.794 24.714 ;
        RECT 34.82 24.672 51.748 24.76 ;
        RECT 43.376 16.116 60.339 16.169 ;
        RECT 51.702 7.79 51.748 24.76 ;
        RECT 34.774 24.718 51.702 24.806 ;
        RECT 43.422 16.07 60.385 16.123 ;
        RECT 51.656 7.836 51.702 24.806 ;
        RECT 34.728 24.764 51.656 24.852 ;
        RECT 43.468 16.024 60.431 16.077 ;
        RECT 51.61 7.882 51.656 24.852 ;
        RECT 34.682 24.81 51.61 24.898 ;
        RECT 43.514 15.978 60.477 16.031 ;
        RECT 51.564 7.928 51.61 24.898 ;
        RECT 34.636 24.856 51.564 24.944 ;
        RECT 43.56 15.932 60.523 15.985 ;
        RECT 51.518 7.974 51.564 24.944 ;
        RECT 34.59 24.902 51.518 24.99 ;
        RECT 43.606 15.886 60.569 15.939 ;
        RECT 51.472 8.02 51.518 24.99 ;
        RECT 34.544 24.948 51.472 25.036 ;
        RECT 43.652 15.84 60.615 15.893 ;
        RECT 51.426 8.066 51.472 25.036 ;
        RECT 34.498 24.994 51.426 25.082 ;
        RECT 43.698 15.794 60.661 15.847 ;
        RECT 51.38 8.112 51.426 25.082 ;
        RECT 34.452 25.04 51.38 25.128 ;
        RECT 43.744 15.748 60.707 15.801 ;
        RECT 51.334 8.158 51.38 25.128 ;
        RECT 34.406 25.086 51.334 25.174 ;
        RECT 43.79 15.702 60.753 15.755 ;
        RECT 51.288 8.204 51.334 25.174 ;
        RECT 34.36 25.132 51.288 25.22 ;
        RECT 43.836 15.656 60.799 15.709 ;
        RECT 51.242 8.25 51.288 25.22 ;
        RECT 34.314 25.178 51.242 25.266 ;
        RECT 43.882 15.61 60.845 15.663 ;
        RECT 51.196 8.296 51.242 25.266 ;
        RECT 34.268 25.224 51.196 25.312 ;
        RECT 43.928 15.564 60.891 15.617 ;
        RECT 51.15 8.342 51.196 25.312 ;
        RECT 34.222 25.27 51.15 25.358 ;
        RECT 43.974 15.518 60.937 15.571 ;
        RECT 51.104 8.388 51.15 25.358 ;
        RECT 34.176 25.316 51.104 25.404 ;
        RECT 44.02 15.472 60.983 15.524 ;
        RECT 51.058 8.434 51.104 25.404 ;
        RECT 34.13 25.362 51.058 25.45 ;
        RECT 44.066 15.426 110 15.5 ;
        RECT 51.012 8.48 51.058 25.45 ;
        RECT 34.084 25.408 51.012 25.496 ;
        RECT 44.112 15.38 110 15.5 ;
        RECT 50.966 8.526 51.012 25.496 ;
        RECT 34.038 25.454 50.966 25.542 ;
        RECT 44.158 15.334 110 15.5 ;
        RECT 50.92 8.572 50.966 25.542 ;
        RECT 33.992 25.5 50.92 25.588 ;
        RECT 44.204 15.288 110 15.5 ;
        RECT 50.874 8.618 50.92 25.588 ;
        RECT 33.946 25.546 50.874 25.634 ;
        RECT 44.25 15.242 110 15.5 ;
        RECT 50.828 8.664 50.874 25.634 ;
        RECT 33.9 25.592 50.828 25.68 ;
        RECT 44.296 15.196 110 15.5 ;
        RECT 50.782 8.71 50.828 25.68 ;
        RECT 33.854 25.638 50.782 25.726 ;
        RECT 44.342 15.15 110 15.5 ;
        RECT 50.736 8.756 50.782 25.726 ;
        RECT 33.808 25.684 50.736 25.772 ;
        RECT 44.388 15.104 110 15.5 ;
        RECT 50.69 8.802 50.736 25.772 ;
        RECT 33.762 25.73 50.69 25.818 ;
        RECT 44.434 15.058 110 15.5 ;
        RECT 50.644 8.848 50.69 25.818 ;
        RECT 33.716 25.776 50.644 25.864 ;
        RECT 44.48 15.012 110 15.5 ;
        RECT 50.598 8.894 50.644 25.864 ;
        RECT 33.67 25.822 50.598 25.91 ;
        RECT 44.526 14.966 110 15.5 ;
        RECT 50.552 8.94 50.598 25.91 ;
        RECT 33.624 25.868 50.552 25.956 ;
        RECT 44.572 14.92 110 15.5 ;
        RECT 50.506 8.986 50.552 25.956 ;
        RECT 33.578 25.914 50.506 26.002 ;
        RECT 44.618 14.874 110 15.5 ;
        RECT 50.46 9.032 50.506 26.002 ;
        RECT 33.532 25.96 50.46 26.048 ;
        RECT 44.664 14.828 110 15.5 ;
        RECT 50.414 9.078 50.46 26.048 ;
        RECT 33.486 26.006 50.414 26.094 ;
        RECT 44.71 14.782 110 15.5 ;
        RECT 50.368 9.124 50.414 26.094 ;
        RECT 33.44 26.052 50.368 26.14 ;
        RECT 44.756 14.736 110 15.5 ;
        RECT 50.322 9.17 50.368 26.14 ;
        RECT 33.394 26.098 50.322 26.186 ;
        RECT 44.802 14.69 110 15.5 ;
        RECT 50.276 9.216 50.322 26.186 ;
        RECT 33.348 26.144 50.276 26.232 ;
        RECT 44.848 14.644 110 15.5 ;
        RECT 50.23 9.262 50.276 26.232 ;
        RECT 33.302 26.19 50.23 26.278 ;
        RECT 44.894 14.598 110 15.5 ;
        RECT 50.184 9.308 50.23 26.278 ;
        RECT 33.256 26.236 50.184 26.324 ;
        RECT 44.94 14.552 110 15.5 ;
        RECT 50.138 9.354 50.184 26.324 ;
        RECT 33.21 26.282 50.138 26.37 ;
        RECT 44.986 14.506 110 15.5 ;
        RECT 50.092 9.4 50.138 26.37 ;
        RECT 33.164 26.328 50.092 26.416 ;
        RECT 45.032 14.46 110 15.5 ;
        RECT 50.046 9.446 50.092 26.416 ;
        RECT 33.118 26.374 50.046 26.462 ;
        RECT 45.078 14.414 110 15.5 ;
        RECT 50 9.492 50.046 26.462 ;
        RECT 33.072 26.42 50 26.508 ;
        RECT 45.124 14.368 110 15.5 ;
        RECT 49.954 9.538 50 26.508 ;
        RECT 33.026 26.466 49.954 26.554 ;
        RECT 45.17 14.322 110 15.5 ;
        RECT 49.908 9.584 49.954 26.554 ;
        RECT 32.98 26.512 49.908 26.6 ;
        RECT 45.216 14.276 110 15.5 ;
        RECT 49.862 9.63 49.908 26.6 ;
        RECT 32.934 26.558 49.862 26.646 ;
        RECT 45.262 14.23 110 15.5 ;
        RECT 49.816 9.676 49.862 26.646 ;
        RECT 32.888 26.604 49.816 26.692 ;
        RECT 45.308 14.184 110 15.5 ;
        RECT 49.77 9.722 49.816 26.692 ;
        RECT 32.842 26.65 49.77 26.738 ;
        RECT 45.354 14.138 110 15.5 ;
        RECT 49.724 9.768 49.77 26.738 ;
        RECT 32.796 26.696 49.724 26.784 ;
        RECT 45.4 14.092 110 15.5 ;
        RECT 49.678 9.814 49.724 26.784 ;
        RECT 32.75 26.742 49.678 26.83 ;
        RECT 45.446 14.046 110 15.5 ;
        RECT 49.632 9.86 49.678 26.83 ;
        RECT 32.704 26.788 49.632 26.876 ;
        RECT 45.492 14 110 15.5 ;
        RECT 49.586 9.906 49.632 26.876 ;
        RECT 32.658 26.834 49.586 26.922 ;
        RECT 45.538 13.954 110 15.5 ;
        RECT 49.54 9.952 49.586 26.922 ;
        RECT 32.612 26.88 49.54 26.968 ;
        RECT 45.584 13.908 110 15.5 ;
        RECT 49.494 9.998 49.54 26.968 ;
        RECT 32.566 26.926 49.494 27.014 ;
        RECT 45.63 13.862 110 15.5 ;
        RECT 49.448 10.044 49.494 27.014 ;
        RECT 32.52 26.972 49.448 27.06 ;
        RECT 45.676 13.816 110 15.5 ;
        RECT 49.402 10.09 49.448 27.06 ;
        RECT 32.474 27.018 49.402 27.106 ;
        RECT 45.722 13.77 110 15.5 ;
        RECT 49.356 10.136 49.402 27.106 ;
        RECT 32.428 27.064 49.356 27.152 ;
        RECT 45.768 13.724 110 15.5 ;
        RECT 49.31 10.182 49.356 27.152 ;
        RECT 32.382 27.11 49.31 27.198 ;
        RECT 45.814 13.678 110 15.5 ;
        RECT 49.264 10.228 49.31 27.198 ;
        RECT 32.336 27.156 49.264 27.244 ;
        RECT 45.86 13.632 110 15.5 ;
        RECT 49.218 10.274 49.264 27.244 ;
        RECT 32.29 27.202 49.218 27.29 ;
        RECT 45.906 13.586 110 15.5 ;
        RECT 49.172 10.32 49.218 27.29 ;
        RECT 32.244 27.248 49.172 27.336 ;
        RECT 45.952 13.54 110 15.5 ;
        RECT 49.126 10.366 49.172 27.336 ;
        RECT 32.198 27.294 49.126 27.382 ;
        RECT 45.998 13.494 110 15.5 ;
        RECT 49.08 10.412 49.126 27.382 ;
        RECT 32.152 27.34 49.08 27.428 ;
        RECT 46.044 13.448 110 15.5 ;
        RECT 49.034 10.458 49.08 27.428 ;
        RECT 32.106 27.386 49.034 27.474 ;
        RECT 46.09 13.402 110 15.5 ;
        RECT 48.988 10.504 49.034 27.474 ;
        RECT 32.06 27.432 48.988 27.52 ;
        RECT 46.136 13.356 110 15.5 ;
        RECT 48.942 10.55 48.988 27.52 ;
        RECT 32.014 27.478 48.942 27.566 ;
        RECT 46.182 13.31 110 15.5 ;
        RECT 48.896 10.596 48.942 27.566 ;
        RECT 31.968 27.524 48.896 27.612 ;
        RECT 46.228 13.264 110 15.5 ;
        RECT 48.85 10.642 48.896 27.612 ;
        RECT 31.922 27.57 48.85 27.658 ;
        RECT 46.274 13.218 110 15.5 ;
        RECT 48.804 10.688 48.85 27.658 ;
        RECT 31.876 27.616 48.804 27.704 ;
        RECT 46.32 13.172 110 15.5 ;
        RECT 48.758 10.734 48.804 27.704 ;
        RECT 31.83 27.662 48.758 27.75 ;
        RECT 46.366 13.126 110 15.5 ;
        RECT 48.712 10.78 48.758 27.75 ;
        RECT 31.784 27.708 48.712 27.796 ;
        RECT 46.412 13.08 110 15.5 ;
        RECT 48.666 10.826 48.712 27.796 ;
        RECT 31.738 27.754 48.666 27.842 ;
        RECT 46.458 13.034 110 15.5 ;
        RECT 48.62 10.872 48.666 27.842 ;
        RECT 31.692 27.8 48.62 27.888 ;
        RECT 46.504 12.988 110 15.5 ;
        RECT 48.574 10.918 48.62 27.888 ;
        RECT 31.646 27.846 48.574 27.934 ;
        RECT 46.55 12.942 110 15.5 ;
        RECT 48.528 10.964 48.574 27.934 ;
        RECT 31.6 27.892 48.528 27.98 ;
        RECT 46.596 12.896 110 15.5 ;
        RECT 48.482 11.01 48.528 27.98 ;
        RECT 31.554 27.938 48.482 28.026 ;
        RECT 46.642 12.85 110 15.5 ;
        RECT 48.436 11.056 48.482 28.026 ;
        RECT 31.508 27.984 48.436 28.072 ;
        RECT 46.688 12.804 110 15.5 ;
        RECT 48.39 11.102 48.436 28.072 ;
        RECT 31.462 28.03 48.39 28.118 ;
        RECT 46.734 12.758 110 15.5 ;
        RECT 48.344 11.148 48.39 28.118 ;
        RECT 31.416 28.076 48.344 28.164 ;
        RECT 46.78 12.712 110 15.5 ;
        RECT 48.298 11.194 48.344 28.164 ;
        RECT 31.37 28.122 48.298 28.21 ;
        RECT 46.826 12.666 110 15.5 ;
        RECT 48.252 11.24 48.298 28.21 ;
        RECT 31.324 28.168 48.252 28.256 ;
        RECT 46.872 12.62 110 15.5 ;
        RECT 48.206 11.286 48.252 28.256 ;
        RECT 31.278 28.214 48.206 28.302 ;
        RECT 46.918 12.574 110 15.5 ;
        RECT 48.16 11.332 48.206 28.302 ;
        RECT 31.232 28.26 48.16 28.348 ;
        RECT 46.964 12.528 110 15.5 ;
        RECT 48.114 11.378 48.16 28.348 ;
        RECT 31.186 28.306 48.114 28.394 ;
        RECT 47.01 12.482 110 15.5 ;
        RECT 48.068 11.424 48.114 28.394 ;
        RECT 31.14 28.352 48.068 28.44 ;
        RECT 47.056 12.436 110 15.5 ;
        RECT 48.022 11.47 48.068 28.44 ;
        RECT 31.094 28.398 48.022 28.486 ;
        RECT 47.102 12.39 110 15.5 ;
        RECT 47.976 11.516 48.022 28.486 ;
        RECT 31.048 28.444 47.976 28.532 ;
        RECT 47.148 12.344 110 15.5 ;
        RECT 47.93 11.562 47.976 28.532 ;
        RECT 31.002 28.49 47.93 28.578 ;
        RECT 47.194 12.298 110 15.5 ;
        RECT 47.884 11.608 47.93 28.578 ;
        RECT 30.956 28.536 47.884 28.624 ;
        RECT 47.24 12.252 110 15.5 ;
        RECT 47.838 11.654 47.884 28.624 ;
        RECT 30.91 28.582 47.838 28.67 ;
        RECT 47.286 12.206 110 15.5 ;
        RECT 47.792 11.7 47.838 28.67 ;
        RECT 30.864 28.628 47.792 28.716 ;
        RECT 47.332 12.16 110 15.5 ;
        RECT 47.746 11.746 47.792 28.716 ;
        RECT 30.818 28.674 47.746 28.762 ;
        RECT 47.378 12.114 110 15.5 ;
        RECT 47.7 11.792 47.746 28.762 ;
        RECT 30.772 28.72 47.7 28.808 ;
        RECT 47.424 12.068 110 15.5 ;
        RECT 47.654 11.838 47.7 28.808 ;
        RECT 30.726 28.766 47.654 28.854 ;
        RECT 47.47 12.022 110 15.5 ;
        RECT 47.608 11.884 47.654 28.854 ;
        RECT 30.68 28.812 47.608 28.9 ;
        RECT 47.516 11.976 110 15.5 ;
        RECT 47.562 11.93 47.608 28.9 ;
        RECT 30.634 28.858 47.562 28.946 ;
        RECT 30.588 28.904 47.516 28.992 ;
        RECT 30.542 28.95 47.47 29.038 ;
        RECT 30.496 28.996 47.424 29.084 ;
        RECT 30.45 29.042 47.378 29.13 ;
        RECT 30.404 29.088 47.332 29.176 ;
        RECT 30.358 29.134 47.286 29.222 ;
        RECT 30.312 29.18 47.24 29.268 ;
        RECT 30.266 29.226 47.194 29.314 ;
        RECT 30.22 29.272 47.148 29.36 ;
        RECT 30.174 29.318 47.102 29.406 ;
        RECT 30.128 29.364 47.056 29.452 ;
        RECT 30.082 29.41 47.01 29.498 ;
        RECT 30.036 29.456 46.964 29.544 ;
        RECT 29.99 29.502 46.918 29.59 ;
        RECT 29.944 29.548 46.872 29.636 ;
        RECT 29.898 29.594 46.826 29.682 ;
        RECT 29.852 29.64 46.78 29.728 ;
        RECT 29.806 29.686 46.734 29.774 ;
        RECT 29.76 29.732 46.688 29.82 ;
        RECT 29.714 29.778 46.642 29.866 ;
        RECT 29.668 29.824 46.596 29.912 ;
        RECT 29.622 29.87 46.55 29.958 ;
        RECT 29.576 29.916 46.504 30.004 ;
        RECT 29.53 29.962 46.458 30.05 ;
        RECT 29.484 30.008 46.412 30.096 ;
        RECT 29.438 30.054 46.366 30.142 ;
        RECT 29.392 30.1 46.32 30.188 ;
        RECT 29.346 30.146 46.274 30.234 ;
        RECT 29.3 30.192 46.228 30.28 ;
        RECT 29.254 30.238 46.182 30.326 ;
        RECT 29.208 30.284 46.136 30.372 ;
        RECT 29.162 30.33 46.09 30.418 ;
        RECT 29.116 30.376 46.044 30.464 ;
        RECT 29.07 30.422 45.998 30.51 ;
        RECT 29.024 30.468 45.952 30.556 ;
        RECT 28.978 30.514 45.906 30.602 ;
        RECT 28.932 30.56 45.86 30.648 ;
        RECT 28.886 30.606 45.814 30.694 ;
        RECT 28.84 30.652 45.768 30.74 ;
        RECT 28.794 30.698 45.722 30.786 ;
        RECT 28.748 30.744 45.676 30.832 ;
        RECT 28.702 30.79 45.63 30.878 ;
        RECT 28.656 30.836 45.584 30.924 ;
        RECT 28.61 30.882 45.538 30.97 ;
        RECT 28.564 30.928 45.492 31.016 ;
        RECT 28.518 30.974 45.446 31.062 ;
        RECT 28.472 31.02 45.4 31.108 ;
        RECT 28.426 31.066 45.354 31.154 ;
        RECT 28.38 31.112 45.308 31.2 ;
        RECT 28.334 31.158 45.262 31.246 ;
        RECT 28.288 31.204 45.216 31.292 ;
        RECT 28.242 31.25 45.17 31.338 ;
        RECT 28.196 31.296 45.124 31.384 ;
        RECT 28.15 31.342 45.078 31.43 ;
        RECT 28.104 31.388 45.032 31.476 ;
        RECT 28.058 31.434 44.986 31.522 ;
        RECT 28.012 31.48 44.94 31.568 ;
        RECT 27.966 31.526 44.894 31.614 ;
        RECT 27.92 31.572 44.848 31.66 ;
        RECT 27.874 31.618 44.802 31.706 ;
        RECT 27.828 31.664 44.756 31.752 ;
        RECT 27.782 31.71 44.71 31.798 ;
        RECT 27.736 31.756 44.664 31.844 ;
        RECT 27.69 31.802 44.618 31.89 ;
        RECT 27.644 31.848 44.572 31.936 ;
        RECT 27.598 31.894 44.526 31.982 ;
        RECT 27.552 31.94 44.48 32.028 ;
        RECT 27.506 31.986 44.434 32.074 ;
        RECT 27.46 32.032 44.388 32.12 ;
        RECT 27.414 32.078 44.342 32.166 ;
        RECT 27.368 32.124 44.296 32.212 ;
        RECT 27.322 32.17 44.25 32.258 ;
        RECT 27.276 32.216 44.204 32.304 ;
        RECT 27.23 32.262 44.158 32.35 ;
        RECT 27.184 32.308 44.112 32.396 ;
        RECT 27.138 32.354 44.066 32.442 ;
        RECT 27.092 32.4 44.02 32.488 ;
        RECT 27.046 32.446 43.974 32.534 ;
        RECT 27 32.492 43.928 32.58 ;
        RECT 26.954 32.538 43.882 32.626 ;
        RECT 26.908 32.584 43.836 32.672 ;
        RECT 26.862 32.63 43.79 32.718 ;
        RECT 26.816 32.676 43.744 32.764 ;
        RECT 26.77 32.722 43.698 32.81 ;
        RECT 26.724 32.768 43.652 32.856 ;
        RECT 26.678 32.814 43.606 32.902 ;
        RECT 26.632 32.86 43.56 32.948 ;
        RECT 26.586 32.906 43.514 32.994 ;
        RECT 26.54 32.952 43.468 33.04 ;
        RECT 26.494 32.998 43.422 33.086 ;
        RECT 26.448 33.044 43.376 33.132 ;
        RECT 26.402 33.09 43.33 33.178 ;
        RECT 26.356 33.136 43.284 33.224 ;
        RECT 26.31 33.182 43.238 33.27 ;
        RECT 26.264 33.228 43.192 33.316 ;
        RECT 26.218 33.274 43.146 33.362 ;
        RECT 26.172 33.32 43.1 33.408 ;
        RECT 26.126 33.366 43.054 33.454 ;
        RECT 26.08 33.412 43.008 33.5 ;
        RECT 26.034 33.458 42.962 33.546 ;
        RECT 25.988 33.504 42.916 33.592 ;
        RECT 25.942 33.55 42.87 33.638 ;
        RECT 25.896 33.596 42.824 33.684 ;
        RECT 25.85 33.642 42.778 33.73 ;
        RECT 25.804 33.688 42.732 33.776 ;
        RECT 25.758 33.734 42.686 33.822 ;
        RECT 25.712 33.78 42.64 33.868 ;
        RECT 25.666 33.826 42.594 33.914 ;
        RECT 25.62 33.872 42.548 33.96 ;
        RECT 25.574 33.918 42.502 34.006 ;
        RECT 25.528 33.964 42.456 34.052 ;
        RECT 25.482 34.01 42.41 34.098 ;
        RECT 25.436 34.056 42.364 34.144 ;
        RECT 25.39 34.102 42.318 34.19 ;
        RECT 25.344 34.148 42.272 34.236 ;
        RECT 25.298 34.194 42.226 34.282 ;
        RECT 25.252 34.24 42.18 34.328 ;
        RECT 25.206 34.286 42.134 34.374 ;
        RECT 25.16 34.332 42.088 34.42 ;
        RECT 25.114 34.378 42.042 34.466 ;
        RECT 25.068 34.424 41.996 34.512 ;
        RECT 25.022 34.47 41.95 34.558 ;
        RECT 24.976 34.516 41.904 34.604 ;
        RECT 24.93 34.562 41.858 34.65 ;
        RECT 24.884 34.608 41.812 34.696 ;
        RECT 24.838 34.654 41.766 34.742 ;
        RECT 24.792 34.7 41.72 34.788 ;
        RECT 24.746 34.746 41.674 34.834 ;
        RECT 24.7 34.792 41.628 34.88 ;
        RECT 24.654 34.838 41.582 34.926 ;
        RECT 24.608 34.884 41.536 34.972 ;
        RECT 24.562 34.93 41.49 35.018 ;
        RECT 24.516 34.976 41.444 35.064 ;
        RECT 24.47 35.022 41.398 35.11 ;
        RECT 24.424 35.068 41.352 35.156 ;
        RECT 24.378 35.114 41.306 35.202 ;
        RECT 24.332 35.16 41.26 35.248 ;
        RECT 24.286 35.206 41.214 35.294 ;
        RECT 24.24 35.252 41.168 35.34 ;
        RECT 24.194 35.298 41.122 35.386 ;
        RECT 24.148 35.344 41.076 35.432 ;
        RECT 24.102 35.39 41.03 35.478 ;
        RECT 24.056 35.436 40.984 35.524 ;
        RECT 24.01 35.482 40.938 35.57 ;
        RECT 23.964 35.528 40.892 35.616 ;
        RECT 23.918 35.574 40.846 35.662 ;
        RECT 23.872 35.62 40.8 35.708 ;
        RECT 23.826 35.666 40.754 35.754 ;
        RECT 23.78 35.712 40.708 35.8 ;
        RECT 23.734 35.758 40.662 35.846 ;
        RECT 23.688 35.804 40.616 35.892 ;
        RECT 23.642 35.85 40.57 35.938 ;
        RECT 23.596 35.896 40.524 35.984 ;
        RECT 23.55 35.942 40.478 36.03 ;
        RECT 23.504 35.988 40.432 36.076 ;
        RECT 23.458 36.034 40.386 36.122 ;
        RECT 23.412 36.08 40.34 36.168 ;
        RECT 23.366 36.126 40.294 36.214 ;
        RECT 23.32 36.172 40.248 36.26 ;
        RECT 23.274 36.218 40.202 36.306 ;
        RECT 23.228 36.264 40.156 36.352 ;
        RECT 23.182 36.31 40.11 36.398 ;
        RECT 23.136 36.356 40.064 36.444 ;
        RECT 23.09 36.402 40.018 36.49 ;
        RECT 23.044 36.448 39.972 36.536 ;
        RECT 22.998 36.494 39.926 36.582 ;
        RECT 22.952 36.54 39.88 36.628 ;
        RECT 22.906 36.586 39.834 36.674 ;
        RECT 22.86 36.632 39.788 36.72 ;
        RECT 22.814 36.678 39.742 36.766 ;
        RECT 22.768 36.724 39.696 36.812 ;
        RECT 22.722 36.77 39.65 36.858 ;
        RECT 22.676 36.816 39.604 36.904 ;
        RECT 22.63 36.862 39.558 36.95 ;
        RECT 22.584 36.908 39.512 36.996 ;
        RECT 22.538 36.954 39.466 37.042 ;
        RECT 22.492 37 39.42 37.088 ;
        RECT 22.446 37.046 39.374 37.134 ;
        RECT 22.4 37.092 39.328 37.18 ;
        RECT 22.354 37.138 39.282 37.226 ;
        RECT 22.308 37.184 39.236 37.272 ;
        RECT 22.262 37.23 39.19 37.318 ;
        RECT 22.216 37.276 39.144 37.364 ;
        RECT 22.17 37.322 39.098 37.41 ;
        RECT 22.124 37.368 39.052 37.456 ;
        RECT 22.078 37.414 39.006 37.502 ;
        RECT 22.032 37.46 38.96 37.548 ;
        RECT 21.986 37.506 38.914 37.594 ;
        RECT 21.94 37.552 38.868 37.64 ;
        RECT 21.894 37.598 38.822 37.686 ;
        RECT 21.848 37.644 38.776 37.732 ;
        RECT 21.802 37.69 38.73 37.778 ;
        RECT 21.756 37.736 38.684 37.824 ;
        RECT 21.71 37.782 38.638 37.87 ;
        RECT 21.664 37.828 38.592 37.916 ;
        RECT 21.618 37.874 38.546 37.962 ;
        RECT 21.572 37.92 38.5 38.008 ;
        RECT 21.526 37.966 38.454 38.054 ;
        RECT 21.48 38.012 38.408 38.1 ;
        RECT 21.434 38.058 38.362 38.146 ;
        RECT 21.388 38.104 38.316 38.192 ;
        RECT 21.342 38.15 38.27 38.238 ;
        RECT 21.296 38.196 38.224 38.284 ;
        RECT 21.25 38.242 38.178 38.33 ;
        RECT 21.204 38.288 38.132 38.376 ;
        RECT 21.158 38.334 38.086 38.422 ;
        RECT 21.112 38.38 38.04 38.468 ;
        RECT 21.066 38.426 37.994 38.514 ;
        RECT 21.02 38.472 37.948 38.56 ;
        RECT 20.974 38.518 37.902 38.606 ;
        RECT 20.928 38.564 37.856 38.652 ;
        RECT 20.882 38.61 37.81 38.698 ;
        RECT 20.836 38.656 37.764 38.744 ;
        RECT 20.79 38.702 37.718 38.79 ;
        RECT 20.744 38.748 37.672 38.836 ;
        RECT 20.698 38.794 37.626 38.882 ;
        RECT 20.652 38.84 37.58 38.928 ;
        RECT 20.606 38.886 37.534 38.974 ;
        RECT 20.56 38.932 37.488 39.02 ;
        RECT 20.514 38.978 37.442 39.066 ;
        RECT 20.468 39.024 37.396 39.112 ;
        RECT 20.422 39.07 37.35 39.158 ;
        RECT 20.376 39.116 37.304 39.204 ;
        RECT 20.33 39.162 37.258 39.25 ;
        RECT 20.284 39.208 37.212 39.296 ;
        RECT 20.238 39.254 37.166 39.342 ;
        RECT 20.192 39.3 37.12 39.388 ;
        RECT 20.146 39.346 37.074 39.434 ;
        RECT 20.1 39.392 37.028 39.48 ;
        RECT 20.054 39.438 36.982 39.526 ;
        RECT 20.008 39.484 36.936 39.572 ;
        RECT 19.962 39.53 36.89 39.618 ;
        RECT 19.916 39.576 36.844 39.664 ;
        RECT 19.87 39.622 36.798 39.71 ;
        RECT 19.824 39.668 36.752 39.756 ;
        RECT 19.778 39.714 36.706 39.802 ;
        RECT 19.732 39.76 36.66 39.848 ;
        RECT 19.686 39.806 36.614 39.894 ;
        RECT 19.64 39.852 36.568 39.94 ;
        RECT 19.594 39.898 36.522 39.986 ;
        RECT 19.548 39.944 36.476 40.032 ;
        RECT 19.502 39.99 36.43 40.078 ;
        RECT 19.456 40.036 36.384 40.124 ;
        RECT 19.41 40.082 36.338 40.17 ;
        RECT 19.364 40.128 36.292 40.216 ;
        RECT 19.318 40.174 36.246 40.262 ;
        RECT 19.272 40.22 36.2 40.308 ;
        RECT 19.226 40.266 36.154 40.354 ;
        RECT 19.18 40.312 36.108 40.4 ;
        RECT 19.134 40.358 36.062 40.446 ;
        RECT 19.088 40.404 36.016 40.492 ;
        RECT 19.042 40.45 35.97 40.538 ;
        RECT 18.996 40.496 35.924 40.584 ;
        RECT 18.95 40.542 35.878 40.63 ;
        RECT 18.904 40.588 35.832 40.676 ;
        RECT 18.858 40.634 35.786 40.722 ;
        RECT 18.812 40.68 35.74 40.768 ;
        RECT 18.766 40.726 35.694 40.814 ;
        RECT 18.72 40.772 35.648 40.86 ;
        RECT 18.674 40.818 35.602 40.906 ;
        RECT 18.628 40.864 35.556 40.952 ;
        RECT 18.582 40.91 35.51 40.998 ;
        RECT 18.536 40.956 35.464 41.044 ;
        RECT 18.49 41.002 35.418 41.09 ;
        RECT 18.444 41.048 35.372 41.136 ;
        RECT 18.398 41.094 35.326 41.182 ;
        RECT 18.352 41.14 35.28 41.228 ;
        RECT 18.306 41.186 35.234 41.274 ;
        RECT 18.26 41.232 35.188 41.32 ;
        RECT 18.214 41.278 35.142 41.366 ;
        RECT 18.168 41.324 35.096 41.412 ;
        RECT 18.122 41.37 35.05 41.458 ;
        RECT 18.076 41.416 35.004 41.504 ;
        RECT 18.03 41.462 34.958 41.55 ;
        RECT 17.984 41.508 34.912 41.596 ;
        RECT 17.938 41.554 34.866 41.642 ;
        RECT 17.892 41.6 34.82 41.688 ;
        RECT 17.846 41.646 34.774 41.734 ;
        RECT 17.8 41.692 34.728 41.78 ;
        RECT 17.754 41.738 34.682 41.826 ;
        RECT 17.708 41.784 34.636 41.872 ;
        RECT 17.662 41.83 34.59 41.918 ;
        RECT 17.616 41.876 34.544 41.964 ;
        RECT 17.57 41.922 34.498 42.01 ;
        RECT 17.524 41.968 34.452 42.056 ;
        RECT 17.478 42.014 34.406 42.102 ;
        RECT 17.432 42.06 34.36 42.148 ;
        RECT 17.386 42.106 34.314 42.194 ;
        RECT 17.34 42.152 34.268 42.24 ;
        RECT 17.294 42.198 34.222 42.286 ;
        RECT 17.248 42.244 34.176 42.332 ;
        RECT 17.202 42.29 34.13 42.378 ;
        RECT 17.156 42.336 34.084 42.424 ;
        RECT 17.11 42.382 34.038 42.47 ;
        RECT 17.064 42.428 33.992 42.516 ;
        RECT 17.018 42.474 33.946 42.562 ;
        RECT 16.972 42.52 33.9 42.608 ;
        RECT 16.926 42.566 33.854 42.654 ;
        RECT 16.88 42.612 33.808 42.7 ;
        RECT 16.834 42.658 33.762 42.746 ;
        RECT 16.788 42.704 33.716 42.792 ;
        RECT 16.742 42.75 33.67 42.838 ;
        RECT 16.696 42.796 33.624 42.884 ;
        RECT 16.65 42.842 33.578 42.93 ;
        RECT 16.604 42.888 33.532 42.976 ;
        RECT 16.558 42.934 33.486 43.022 ;
        RECT 16.512 42.98 33.44 43.068 ;
        RECT 16.466 43.026 33.394 43.114 ;
        RECT 16.42 43.072 33.348 43.16 ;
        RECT 16.374 43.118 33.302 43.206 ;
        RECT 16.328 43.164 33.256 43.252 ;
        RECT 16.282 43.21 33.21 43.298 ;
        RECT 16.236 43.256 33.164 43.344 ;
        RECT 16.19 43.302 33.118 43.39 ;
        RECT 16.144 43.348 33.072 43.436 ;
        RECT 16.098 43.394 33.026 43.482 ;
        RECT 16.052 43.44 32.98 43.528 ;
        RECT 16.006 43.486 32.934 43.574 ;
        RECT 15.96 43.532 32.888 43.62 ;
        RECT 15.914 43.578 32.842 43.666 ;
        RECT 15.868 43.624 32.796 43.712 ;
        RECT 15.822 43.67 32.75 43.758 ;
        RECT 15.776 43.716 32.704 43.804 ;
        RECT 15.73 43.762 32.658 43.85 ;
        RECT 15.684 43.808 32.612 43.896 ;
        RECT 15.638 43.854 32.566 43.942 ;
        RECT 15.592 43.9 32.52 43.988 ;
        RECT 15.5 43.992 32.474 44.034 ;
        RECT 15.546 43.946 32.474 44.034 ;
        RECT 15.46 44.035 32.428 44.08 ;
        RECT 15.414 44.078 32.382 44.126 ;
        RECT 15.368 44.124 32.336 44.172 ;
        RECT 15.322 44.17 32.29 44.218 ;
        RECT 15.276 44.216 32.244 44.264 ;
        RECT 15.23 44.262 32.198 44.31 ;
        RECT 15.184 44.308 32.152 44.356 ;
        RECT 15.138 44.354 32.106 44.402 ;
        RECT 15.092 44.4 32.06 44.448 ;
        RECT 15.046 44.446 32.014 44.494 ;
        RECT 15 44.492 31.968 44.54 ;
        RECT 14.954 44.538 31.922 44.586 ;
        RECT 14.908 44.584 31.876 44.632 ;
        RECT 14.862 44.63 31.83 44.678 ;
        RECT 14.816 44.676 31.784 44.724 ;
        RECT 14.77 44.722 31.738 44.77 ;
        RECT 14.724 44.768 31.692 44.816 ;
        RECT 14.678 44.814 31.646 44.862 ;
        RECT 14.632 44.86 31.6 44.908 ;
        RECT 14.586 44.906 31.554 44.954 ;
        RECT 14.54 44.952 31.508 45 ;
        RECT 14.494 44.998 31.462 45.046 ;
        RECT 14.448 45.044 31.416 45.092 ;
        RECT 14.402 45.09 31.37 45.138 ;
        RECT 14.356 45.136 31.324 45.184 ;
        RECT 14.31 45.182 31.278 45.23 ;
        RECT 14.264 45.228 31.232 45.276 ;
        RECT 14.218 45.274 31.186 45.322 ;
        RECT 14.172 45.32 31.14 45.368 ;
        RECT 14.126 45.366 31.094 45.414 ;
        RECT 14.08 45.412 31.048 45.46 ;
        RECT 14.034 45.458 31.002 45.506 ;
        RECT 13.988 45.504 30.956 45.552 ;
        RECT 13.942 45.55 30.91 45.598 ;
        RECT 13.896 45.596 30.864 45.644 ;
        RECT 13.85 45.642 30.818 45.69 ;
        RECT 13.804 45.688 30.772 45.736 ;
        RECT 13.758 45.734 30.726 45.782 ;
        RECT 13.712 45.78 30.68 45.828 ;
        RECT 13.666 45.826 30.634 45.874 ;
        RECT 13.62 45.872 30.588 45.92 ;
        RECT 13.574 45.918 30.542 45.966 ;
        RECT 13.528 45.964 30.496 46.012 ;
        RECT 13.482 46.01 30.45 46.058 ;
        RECT 13.436 46.056 30.404 46.104 ;
        RECT 13.39 46.102 30.358 46.15 ;
        RECT 13.344 46.148 30.312 46.196 ;
        RECT 13.298 46.194 30.266 46.242 ;
        RECT 13.252 46.24 30.22 46.288 ;
        RECT 13.206 46.286 30.174 46.334 ;
        RECT 13.16 46.332 30.128 46.38 ;
        RECT 13.114 46.378 30.082 46.426 ;
        RECT 13.068 46.424 30.036 46.472 ;
        RECT 13.022 46.47 29.99 46.518 ;
        RECT 12.976 46.516 29.944 46.564 ;
        RECT 12.93 46.562 29.898 46.61 ;
        RECT 12.884 46.608 29.852 46.656 ;
        RECT 12.838 46.654 29.806 46.702 ;
        RECT 12.792 46.7 29.76 46.748 ;
        RECT 12.746 46.746 29.714 46.794 ;
        RECT 12.7 46.792 29.668 46.84 ;
        RECT 12.654 46.838 29.622 46.886 ;
        RECT 12.608 46.884 29.576 46.932 ;
        RECT 12.562 46.93 29.53 46.978 ;
        RECT 12.516 46.976 29.484 47.024 ;
        RECT 12.47 47.022 29.438 47.07 ;
        RECT 12.424 47.068 29.392 47.116 ;
        RECT 12.378 47.114 29.346 47.162 ;
        RECT 12.332 47.16 29.3 47.208 ;
        RECT 12.286 47.206 29.254 47.254 ;
        RECT 12.24 47.252 29.208 47.3 ;
        RECT 12.194 47.298 29.162 47.346 ;
        RECT 12.148 47.344 29.116 47.392 ;
        RECT 12.102 47.39 29.07 47.438 ;
        RECT 12.056 47.436 29.024 47.484 ;
        RECT 12.01 47.482 28.978 47.53 ;
        RECT 11.964 47.528 28.932 47.576 ;
        RECT 11.918 47.574 28.886 47.622 ;
        RECT 11.872 47.62 28.84 47.668 ;
        RECT 11.826 47.666 28.794 47.714 ;
        RECT 11.78 47.712 28.748 47.76 ;
        RECT 11.734 47.758 28.702 47.806 ;
        RECT 11.688 47.804 28.656 47.852 ;
        RECT 11.642 47.85 28.61 47.898 ;
        RECT 11.596 47.896 28.564 47.944 ;
        RECT 11.55 47.942 28.518 47.99 ;
        RECT 11.504 47.988 28.472 48.036 ;
        RECT 11.458 48.034 28.426 48.082 ;
        RECT 11.412 48.08 28.38 48.128 ;
        RECT 11.366 48.126 28.334 48.174 ;
        RECT 11.32 48.172 28.288 48.22 ;
        RECT 11.274 48.218 28.242 48.266 ;
        RECT 11.228 48.264 28.196 48.312 ;
        RECT 11.182 48.31 28.15 48.358 ;
        RECT 11.136 48.356 28.104 48.404 ;
        RECT 11.09 48.402 28.058 48.45 ;
        RECT 11.044 48.448 28.012 48.496 ;
        RECT 10.998 48.494 27.966 48.542 ;
        RECT 10.952 48.54 27.92 48.588 ;
        RECT 10.906 48.586 27.874 48.634 ;
        RECT 10.86 48.632 27.828 48.68 ;
        RECT 10.814 48.678 27.782 48.726 ;
        RECT 10.768 48.724 27.736 48.772 ;
        RECT 10.722 48.77 27.69 48.818 ;
        RECT 10.676 48.816 27.644 48.864 ;
        RECT 10.63 48.862 27.598 48.91 ;
        RECT 10.584 48.908 27.552 48.956 ;
        RECT 10.538 48.954 27.506 49.002 ;
        RECT 10.492 49 27.46 49.048 ;
        RECT 10.446 49.046 27.414 49.094 ;
        RECT 10.4 49.092 27.368 49.14 ;
        RECT 10.354 49.138 27.322 49.186 ;
        RECT 10.308 49.184 27.276 49.232 ;
        RECT 10.262 49.23 27.23 49.278 ;
        RECT 10.216 49.276 27.184 49.324 ;
        RECT 10.17 49.322 27.138 49.37 ;
        RECT 10.124 49.368 27.092 49.416 ;
        RECT 10.078 49.414 27.046 49.462 ;
      LAYER MET3 ;
        RECT 28.362 51.38 45.33 51.428 ;
        RECT 28.316 51.426 45.284 51.474 ;
        RECT 28.27 51.472 45.238 51.52 ;
        RECT 28.224 51.518 45.192 51.566 ;
        RECT 28.178 51.564 45.146 51.612 ;
        RECT 28.132 51.61 45.1 51.658 ;
        RECT 28.086 51.656 45.054 51.704 ;
        RECT 28.04 51.702 45.008 51.75 ;
        RECT 27.994 51.748 44.962 51.796 ;
        RECT 27.948 51.794 44.916 51.842 ;
        RECT 27.902 51.84 44.87 51.888 ;
        RECT 27.856 51.886 44.824 51.934 ;
        RECT 27.81 51.932 44.778 51.98 ;
        RECT 27.764 51.978 44.732 52.026 ;
        RECT 27.718 52.024 44.686 52.072 ;
        RECT 27.672 52.07 44.64 52.118 ;
        RECT 27.626 52.116 44.594 52.164 ;
        RECT 27.58 52.162 44.548 52.21 ;
        RECT 27.534 52.208 44.502 52.256 ;
        RECT 27.488 52.254 44.456 52.302 ;
        RECT 27.442 52.3 44.41 52.348 ;
        RECT 27.396 52.346 44.364 52.394 ;
        RECT 27.35 52.392 44.318 52.44 ;
        RECT 27.304 52.438 44.272 52.486 ;
        RECT 27.258 52.484 44.226 52.532 ;
        RECT 27.212 52.53 44.18 52.578 ;
        RECT 27.166 52.576 44.134 52.624 ;
        RECT 27.12 52.622 44.088 52.67 ;
        RECT 27.074 52.668 44.042 52.716 ;
        RECT 27.028 52.714 43.996 52.762 ;
        RECT 26.982 52.76 43.95 52.808 ;
        RECT 26.936 52.806 43.904 52.854 ;
        RECT 26.89 52.852 43.858 52.9 ;
        RECT 26.844 52.898 43.812 52.946 ;
        RECT 26.798 52.944 43.766 52.992 ;
        RECT 26.752 52.99 43.72 53.038 ;
        RECT 26.706 53.036 43.674 53.084 ;
        RECT 26.66 53.082 43.628 53.13 ;
        RECT 26.614 53.128 43.582 53.176 ;
        RECT 26.568 53.174 43.536 53.222 ;
        RECT 26.522 53.22 43.49 53.268 ;
        RECT 26.476 53.266 43.444 53.314 ;
        RECT 26.43 53.312 43.398 53.36 ;
        RECT 26.384 53.358 43.352 53.406 ;
        RECT 26.338 53.404 43.306 53.452 ;
        RECT 26.292 53.45 43.26 53.498 ;
        RECT 26.246 53.496 43.214 53.544 ;
        RECT 26.2 53.542 43.168 53.59 ;
        RECT 26.154 53.588 43.122 53.636 ;
        RECT 26.108 53.634 43.076 53.682 ;
        RECT 26.062 53.68 43.03 53.728 ;
        RECT 26.016 53.726 42.984 53.774 ;
        RECT 25.97 53.772 42.938 53.82 ;
        RECT 25.924 53.818 42.892 53.866 ;
        RECT 25.878 53.864 42.846 53.912 ;
        RECT 25.832 53.91 42.8 53.958 ;
        RECT 25.786 53.956 42.754 54.004 ;
        RECT 25.74 54.002 42.708 54.05 ;
        RECT 25.694 54.048 42.662 54.096 ;
        RECT 25.648 54.094 42.616 54.142 ;
        RECT 25.602 54.14 42.57 54.188 ;
        RECT 25.556 54.186 42.524 54.234 ;
        RECT 25.51 54.232 42.478 54.28 ;
        RECT 25.464 54.278 42.432 54.326 ;
        RECT 25.418 54.324 42.386 54.372 ;
        RECT 25.372 54.37 42.34 54.418 ;
        RECT 25.326 54.416 42.294 54.464 ;
        RECT 25.28 54.462 42.248 54.51 ;
        RECT 25.234 54.508 42.202 54.556 ;
        RECT 25.188 54.554 42.156 54.602 ;
        RECT 25.142 54.6 42.11 54.648 ;
        RECT 25.096 54.646 42.064 54.694 ;
        RECT 25.05 54.692 42.018 54.74 ;
        RECT 25.004 54.738 41.972 54.786 ;
        RECT 24.958 54.784 41.926 54.832 ;
        RECT 24.912 54.83 41.88 54.878 ;
        RECT 24.866 54.876 41.834 54.924 ;
        RECT 24.82 54.922 41.788 54.97 ;
        RECT 24.774 54.968 41.742 55.016 ;
        RECT 24.728 55.014 41.696 55.062 ;
        RECT 24.682 55.06 41.65 55.108 ;
        RECT 24.636 55.106 41.604 55.154 ;
        RECT 24.59 55.152 41.558 55.2 ;
        RECT 24.544 55.198 41.512 55.246 ;
        RECT 24.498 55.244 41.466 55.292 ;
        RECT 24.452 55.29 41.42 55.338 ;
        RECT 24.406 55.336 41.374 55.384 ;
        RECT 24.36 55.382 41.328 55.43 ;
        RECT 24.314 55.428 41.282 55.476 ;
        RECT 24.268 55.474 41.236 55.522 ;
        RECT 24.222 55.52 41.19 55.568 ;
        RECT 24.176 55.566 41.144 55.614 ;
        RECT 24.13 55.612 41.098 55.66 ;
        RECT 24.084 55.658 41.052 55.706 ;
        RECT 24.038 55.704 41.006 55.752 ;
        RECT 23.992 55.75 40.96 55.798 ;
        RECT 23.946 55.796 40.914 55.844 ;
        RECT 23.9 55.842 40.868 55.89 ;
        RECT 23.854 55.888 40.822 55.936 ;
        RECT 23.808 55.934 40.776 55.982 ;
        RECT 23.762 55.98 40.73 56.028 ;
        RECT 23.716 56.026 40.684 56.074 ;
        RECT 23.67 56.072 40.638 56.12 ;
        RECT 23.624 56.118 40.592 56.166 ;
        RECT 23.578 56.164 40.546 56.212 ;
        RECT 23.532 56.21 40.5 56.258 ;
        RECT 23.486 56.256 40.454 56.304 ;
        RECT 23.44 56.302 40.408 56.35 ;
        RECT 23.394 56.348 40.362 56.396 ;
        RECT 23.348 56.394 40.316 56.442 ;
        RECT 23.302 56.44 40.27 56.488 ;
        RECT 23.256 56.486 40.224 56.534 ;
        RECT 23.21 56.532 40.178 56.58 ;
        RECT 23.164 56.578 40.132 56.626 ;
        RECT 23.118 56.624 40.086 56.672 ;
        RECT 23.072 56.67 40.04 56.718 ;
        RECT 23.026 56.716 39.994 56.764 ;
        RECT 22.98 56.762 39.948 56.81 ;
        RECT 22.934 56.808 39.902 56.856 ;
        RECT 22.888 56.854 39.856 56.902 ;
        RECT 22.842 56.9 39.81 56.948 ;
        RECT 22.796 56.946 39.764 56.994 ;
        RECT 22.75 56.992 39.718 57.04 ;
        RECT 22.704 57.038 39.672 57.086 ;
        RECT 22.658 57.084 39.626 57.132 ;
        RECT 22.612 57.13 39.58 57.178 ;
        RECT 22.566 57.176 39.534 57.224 ;
        RECT 22.52 57.222 39.488 57.27 ;
        RECT 22.474 57.268 39.442 57.316 ;
        RECT 22.428 57.314 39.396 57.362 ;
        RECT 22.382 57.36 39.35 57.408 ;
        RECT 22.336 57.406 39.304 57.454 ;
        RECT 22.29 57.452 39.258 57.5 ;
        RECT 22.244 57.498 39.212 57.546 ;
        RECT 22.198 57.544 39.166 57.592 ;
        RECT 22.152 57.59 39.12 57.638 ;
        RECT 22.106 57.636 39.074 57.684 ;
        RECT 22.06 57.682 39.028 57.73 ;
        RECT 22.014 57.728 38.982 57.776 ;
        RECT 21.968 57.774 38.936 57.822 ;
        RECT 21.922 57.82 38.89 57.868 ;
        RECT 21.876 57.866 38.844 57.914 ;
        RECT 21.83 57.912 38.798 57.96 ;
        RECT 21.784 57.958 38.752 58.006 ;
        RECT 21.738 58.004 38.706 58.052 ;
        RECT 21.692 58.05 38.66 58.098 ;
        RECT 21.646 58.096 38.614 58.144 ;
        RECT 21.6 58.142 38.568 58.19 ;
        RECT 21.554 58.188 38.522 58.236 ;
        RECT 21.508 58.234 38.476 58.282 ;
        RECT 21.462 58.28 38.43 58.328 ;
        RECT 21.416 58.326 38.384 58.374 ;
        RECT 21.37 58.372 38.338 58.42 ;
        RECT 21.324 58.418 38.292 58.466 ;
        RECT 21.278 58.464 38.246 58.512 ;
        RECT 21.232 58.51 38.2 58.558 ;
        RECT 21.186 58.556 38.154 58.604 ;
        RECT 21.14 58.602 38.108 58.65 ;
        RECT 21.094 58.648 38.062 58.696 ;
        RECT 21.048 58.694 38.016 58.742 ;
        RECT 21.002 58.74 37.97 58.788 ;
        RECT 20.956 58.786 37.924 58.834 ;
        RECT 20.91 58.832 37.878 58.88 ;
        RECT 20.864 58.878 37.832 58.926 ;
        RECT 20.818 58.924 37.786 58.972 ;
        RECT 20.772 58.97 37.74 59.018 ;
        RECT 20.726 59.016 37.694 59.064 ;
        RECT 20.68 59.062 37.648 59.11 ;
        RECT 20.634 59.108 37.602 59.156 ;
        RECT 20.588 59.154 37.556 59.202 ;
        RECT 20.542 59.2 37.51 59.248 ;
        RECT 20.496 59.246 37.464 59.294 ;
        RECT 20.45 59.292 37.418 59.34 ;
        RECT 20.404 59.338 37.372 59.386 ;
        RECT 20.358 59.384 37.326 59.432 ;
        RECT 20.312 59.43 37.28 59.478 ;
        RECT 20.266 59.476 37.234 59.524 ;
        RECT 20.22 59.522 37.188 59.57 ;
        RECT 20.174 59.568 37.142 59.616 ;
        RECT 20.128 59.614 37.096 59.662 ;
        RECT 20.082 59.66 37.05 59.708 ;
        RECT 20.036 59.706 37.004 59.754 ;
        RECT 19.99 59.752 36.958 59.8 ;
        RECT 19.944 59.798 36.912 59.846 ;
        RECT 19.898 59.844 36.866 59.892 ;
        RECT 19.852 59.89 36.82 59.938 ;
        RECT 19.806 59.936 36.774 59.984 ;
        RECT 19.76 59.982 36.728 60.03 ;
        RECT 19.714 60.028 36.682 60.076 ;
        RECT 19.668 60.074 36.636 60.122 ;
        RECT 19.622 60.12 36.59 60.168 ;
        RECT 19.576 60.166 36.544 60.214 ;
        RECT 19.53 60.212 36.498 60.26 ;
        RECT 19.484 60.258 36.452 60.306 ;
        RECT 19.438 60.304 36.406 60.352 ;
        RECT 19.392 60.35 36.36 60.398 ;
        RECT 19.346 60.396 36.314 60.444 ;
        RECT 19.3 60.442 36.268 60.49 ;
        RECT 19.254 60.488 36.222 60.536 ;
        RECT 19.208 60.534 36.176 60.582 ;
        RECT 19.162 60.58 36.13 60.628 ;
        RECT 19.116 60.626 36.084 60.674 ;
        RECT 19.07 60.672 36.038 60.72 ;
        RECT 19.024 60.718 35.992 60.766 ;
        RECT 18.978 60.764 35.946 60.812 ;
        RECT 18.932 60.81 35.9 60.858 ;
        RECT 18.886 60.856 35.854 60.904 ;
        RECT 18.84 60.902 35.808 60.95 ;
        RECT 18.794 60.948 35.762 60.996 ;
        RECT 18.748 60.994 35.716 61.042 ;
        RECT 18.702 61.04 35.67 61.088 ;
        RECT 18.656 61.086 35.624 61.134 ;
        RECT 18.61 61.132 35.578 61.18 ;
        RECT 18.564 61.178 35.532 61.226 ;
        RECT 18.518 61.224 35.486 61.272 ;
        RECT 18.472 61.27 35.44 61.318 ;
        RECT 18.426 61.316 35.394 61.364 ;
        RECT 18.38 61.362 35.348 61.41 ;
        RECT 18.334 61.408 35.302 61.456 ;
        RECT 18.288 61.454 35.256 61.502 ;
        RECT 18.242 61.5 35.21 61.548 ;
        RECT 18.196 61.546 35.164 61.594 ;
        RECT 18.15 61.592 35.118 61.64 ;
        RECT 18.104 61.638 35.072 61.686 ;
        RECT 18.058 61.684 35.026 61.732 ;
        RECT 18.012 61.73 34.98 61.778 ;
        RECT 17.966 61.776 34.934 61.824 ;
        RECT 17.92 61.822 34.888 61.87 ;
        RECT 17.874 61.868 34.842 61.916 ;
        RECT 17.828 61.914 34.796 61.962 ;
        RECT 17.782 61.96 34.75 62.008 ;
        RECT 17.736 62.006 34.704 62.054 ;
        RECT 17.69 62.052 34.658 62.1 ;
        RECT 17.644 62.098 34.612 62.146 ;
        RECT 17.598 62.144 34.566 62.192 ;
        RECT 17.552 62.19 34.52 62.238 ;
        RECT 17.506 62.236 34.474 62.284 ;
        RECT 17.46 62.282 34.428 62.33 ;
        RECT 17.414 62.328 34.382 62.376 ;
        RECT 17.368 62.374 34.336 62.422 ;
        RECT 17.322 62.42 34.29 62.468 ;
        RECT 17.276 62.466 34.244 62.514 ;
        RECT 17.23 62.512 34.198 62.56 ;
        RECT 17.184 62.558 34.152 62.606 ;
        RECT 17.138 62.604 34.106 62.652 ;
        RECT 17.092 62.65 34.06 62.698 ;
        RECT 17.046 62.696 34.014 62.744 ;
        RECT 17 62.742 33.968 62.79 ;
        RECT 17 62.742 33.922 62.836 ;
        RECT 17 62.742 33.876 62.882 ;
        RECT 17 62.742 33.83 62.928 ;
        RECT 17 62.742 33.784 62.974 ;
        RECT 17 62.742 33.738 63.02 ;
        RECT 17 62.742 33.692 63.066 ;
        RECT 17 62.742 33.646 63.112 ;
        RECT 17 62.742 33.6 63.158 ;
        RECT 17 62.742 33.554 63.204 ;
        RECT 17 62.742 33.508 63.25 ;
        RECT 17 62.742 33.462 63.296 ;
        RECT 17 62.742 33.416 63.342 ;
        RECT 17 62.742 33.37 63.388 ;
        RECT 17 62.742 33.324 63.434 ;
        RECT 17 62.742 33.278 63.48 ;
        RECT 17 62.742 33.232 63.526 ;
        RECT 17 62.742 33.186 63.572 ;
        RECT 17 62.742 33.14 63.618 ;
        RECT 17 62.742 33.094 63.664 ;
        RECT 17 62.742 33.048 63.71 ;
        RECT 17 62.742 33.002 63.756 ;
        RECT 17 62.742 32.956 63.802 ;
        RECT 17 62.742 32.91 63.848 ;
        RECT 17 62.742 32.864 63.894 ;
        RECT 17 62.742 32.818 63.94 ;
        RECT 17 62.742 32.772 63.986 ;
        RECT 17 62.742 32.726 64.032 ;
        RECT 17 62.742 32.68 64.078 ;
        RECT 17 62.742 32.634 64.124 ;
        RECT 17 62.742 32.588 64.17 ;
        RECT 17 62.742 32.542 64.216 ;
        RECT 17 62.742 32.496 64.262 ;
        RECT 17 62.742 32.45 64.308 ;
        RECT 17 62.742 32.404 64.354 ;
        RECT 17 62.742 32.358 64.4 ;
        RECT 17 62.742 32.312 64.446 ;
        RECT 17 62.742 32.266 64.492 ;
        RECT 17 62.742 32.22 64.538 ;
        RECT 17 62.742 32.174 64.584 ;
        RECT 17 62.742 32.128 64.63 ;
        RECT 17 62.742 32.082 64.676 ;
        RECT 17 62.742 32.036 64.722 ;
        RECT 17 62.742 31.99 64.768 ;
        RECT 17 62.742 31.944 64.814 ;
        RECT 17 62.742 31.898 64.86 ;
        RECT 17 62.742 31.852 64.906 ;
        RECT 17 62.742 31.806 64.952 ;
        RECT 17 62.742 31.76 64.998 ;
        RECT 17 62.742 31.714 65.044 ;
        RECT 17 62.742 31.668 65.09 ;
        RECT 17 62.742 31.622 65.136 ;
        RECT 17 62.742 31.576 65.182 ;
        RECT 17 62.742 31.53 65.228 ;
        RECT 17 62.742 31.484 65.274 ;
        RECT 17 62.742 31.438 65.32 ;
        RECT 17 62.742 31.392 65.366 ;
        RECT 17 62.742 31.346 65.412 ;
        RECT 17 62.742 31.3 65.458 ;
        RECT 17 62.742 31.254 65.504 ;
        RECT 17 62.742 31.208 65.55 ;
        RECT 17 62.742 31.162 65.596 ;
        RECT 17 62.742 31.116 65.642 ;
        RECT 17 62.742 31.07 65.688 ;
        RECT 17 62.742 31.024 65.734 ;
        RECT 17 62.742 30.978 65.78 ;
        RECT 17 62.742 30.932 65.826 ;
        RECT 17 62.742 30.886 65.872 ;
        RECT 17 62.742 30.84 65.918 ;
        RECT 17 62.742 30.794 65.964 ;
        RECT 17 62.742 30.748 66.01 ;
        RECT 17 62.742 30.702 66.056 ;
        RECT 17 62.742 30.656 66.102 ;
        RECT 17 62.742 30.61 66.148 ;
        RECT 17 62.742 30.564 66.194 ;
        RECT 17 62.742 30.518 66.24 ;
        RECT 17 62.742 30.472 66.286 ;
        RECT 17 62.742 30.426 66.332 ;
        RECT 17 62.742 30.38 66.378 ;
        RECT 17 62.742 30.334 66.424 ;
        RECT 17 62.742 30.288 66.47 ;
        RECT 17 62.742 30.242 66.516 ;
        RECT 17 62.742 30.196 66.562 ;
        RECT 17 62.742 30.15 66.608 ;
        RECT 17 62.742 30.104 66.654 ;
        RECT 17 62.742 30.058 66.7 ;
        RECT 17 62.742 30.012 66.746 ;
        RECT 17 62.742 29.966 66.792 ;
        RECT 17 62.742 29.92 66.838 ;
        RECT 17 62.742 29.874 66.884 ;
        RECT 17 62.742 29.828 66.93 ;
        RECT 17 62.742 29.782 66.976 ;
        RECT 17 62.742 29.736 67.022 ;
        RECT 17 62.742 29.69 67.068 ;
        RECT 17 62.742 29.644 67.114 ;
        RECT 17 62.742 29.598 67.16 ;
        RECT 17 62.742 29.552 67.206 ;
        RECT 17 62.742 29.506 67.252 ;
        RECT 17 62.742 29.46 67.298 ;
        RECT 17 62.742 29.414 67.344 ;
        RECT 17 62.742 29.368 67.39 ;
        RECT 17 62.742 29.322 67.436 ;
        RECT 17 62.742 29.276 67.482 ;
        RECT 17 62.742 29.23 67.528 ;
        RECT 17 62.742 29.184 67.574 ;
        RECT 17 62.742 29.138 67.62 ;
        RECT 17 62.742 29.092 67.666 ;
        RECT 17 62.742 29.046 67.712 ;
        RECT 17 62.742 29 110 ;
        RECT 92.47 78.5 110 89.5 ;
        RECT 81.444 89.503 97.024 89.529 ;
        RECT 78.5 92.447 94.034 92.519 ;
        RECT 78.5 92.447 93.988 92.565 ;
        RECT 78.5 92.447 93.942 92.611 ;
        RECT 78.5 92.447 93.896 92.657 ;
        RECT 78.5 92.447 93.85 92.703 ;
        RECT 78.5 92.447 93.804 92.749 ;
        RECT 78.5 92.447 93.758 92.795 ;
        RECT 78.5 92.447 93.712 92.841 ;
        RECT 78.5 92.447 93.666 92.887 ;
        RECT 78.5 92.447 93.62 92.933 ;
        RECT 78.5 92.447 93.574 92.979 ;
        RECT 78.5 92.447 93.528 93.025 ;
        RECT 78.5 92.447 93.482 93.071 ;
        RECT 78.5 92.447 93.436 93.117 ;
        RECT 78.5 92.447 93.39 93.163 ;
        RECT 78.5 92.447 93.344 93.209 ;
        RECT 78.5 92.447 93.298 93.255 ;
        RECT 78.5 92.447 93.252 93.301 ;
        RECT 78.5 92.447 93.206 93.347 ;
        RECT 78.5 92.447 93.16 93.393 ;
        RECT 78.5 92.447 93.114 93.439 ;
        RECT 78.5 92.447 93.068 93.485 ;
        RECT 78.5 92.447 93.022 93.531 ;
        RECT 78.5 92.447 92.976 93.577 ;
        RECT 78.5 92.447 92.93 93.623 ;
        RECT 78.5 92.447 92.884 93.669 ;
        RECT 78.5 92.447 92.838 93.715 ;
        RECT 78.5 92.447 92.792 93.761 ;
        RECT 78.5 92.447 92.746 93.807 ;
        RECT 78.5 92.447 92.7 93.853 ;
        RECT 78.5 92.447 92.654 93.899 ;
        RECT 78.5 92.447 92.608 93.945 ;
        RECT 78.5 92.447 92.562 93.991 ;
        RECT 78.5 92.447 92.516 94.037 ;
        RECT 78.546 92.401 94.08 92.473 ;
        RECT 92.444 78.513 92.47 94.073 ;
        RECT 78.592 92.355 94.126 92.427 ;
        RECT 92.398 78.549 92.444 94.109 ;
        RECT 78.638 92.309 94.172 92.381 ;
        RECT 92.352 78.595 92.398 94.155 ;
        RECT 78.684 92.263 94.218 92.335 ;
        RECT 92.306 78.641 92.352 94.201 ;
        RECT 78.73 92.217 94.264 92.289 ;
        RECT 92.26 78.687 92.306 94.247 ;
        RECT 78.776 92.171 94.31 92.243 ;
        RECT 92.214 78.733 92.26 94.293 ;
        RECT 78.822 92.125 94.356 92.197 ;
        RECT 92.168 78.779 92.214 94.339 ;
        RECT 78.868 92.079 94.402 92.151 ;
        RECT 92.122 78.825 92.168 94.385 ;
        RECT 78.914 92.033 94.448 92.105 ;
        RECT 92.076 78.871 92.122 94.431 ;
        RECT 78.96 91.987 94.494 92.059 ;
        RECT 92.03 78.917 92.076 94.477 ;
        RECT 79.006 91.941 94.54 92.013 ;
        RECT 91.984 78.963 92.03 94.523 ;
        RECT 79.052 91.895 94.586 91.967 ;
        RECT 91.938 79.009 91.984 94.569 ;
        RECT 79.098 91.849 94.632 91.921 ;
        RECT 91.892 79.055 91.938 94.615 ;
        RECT 79.144 91.803 94.678 91.875 ;
        RECT 91.846 79.101 91.892 94.661 ;
        RECT 79.19 91.757 94.724 91.829 ;
        RECT 91.8 79.147 91.846 94.707 ;
        RECT 79.236 91.711 94.77 91.783 ;
        RECT 91.754 79.193 91.8 94.753 ;
        RECT 79.282 91.665 94.816 91.737 ;
        RECT 91.708 79.239 91.754 94.799 ;
        RECT 79.328 91.619 94.862 91.691 ;
        RECT 91.662 79.285 91.708 94.845 ;
        RECT 79.374 91.573 94.908 91.645 ;
        RECT 91.616 79.331 91.662 94.891 ;
        RECT 79.42 91.527 94.954 91.599 ;
        RECT 91.57 79.377 91.616 94.937 ;
        RECT 79.466 91.481 95 91.553 ;
        RECT 91.524 79.423 91.57 94.983 ;
        RECT 79.512 91.435 95.046 91.507 ;
        RECT 91.478 79.469 91.524 95.029 ;
        RECT 79.558 91.389 95.092 91.461 ;
        RECT 91.432 79.515 91.478 95.075 ;
        RECT 79.604 91.343 95.138 91.415 ;
        RECT 91.386 79.561 91.432 95.121 ;
        RECT 79.65 91.297 95.184 91.369 ;
        RECT 91.34 79.607 91.386 95.167 ;
        RECT 79.696 91.251 95.23 91.323 ;
        RECT 91.294 79.653 91.34 95.213 ;
        RECT 79.742 91.205 95.276 91.277 ;
        RECT 91.248 79.699 91.294 95.259 ;
        RECT 79.788 91.159 95.322 91.231 ;
        RECT 91.202 79.745 91.248 95.305 ;
        RECT 79.834 91.113 95.368 91.185 ;
        RECT 91.156 79.791 91.202 95.351 ;
        RECT 79.88 91.067 95.414 91.139 ;
        RECT 91.11 79.837 91.156 95.397 ;
        RECT 79.926 91.021 95.46 91.093 ;
        RECT 91.064 79.883 91.11 95.443 ;
        RECT 79.972 90.975 95.506 91.047 ;
        RECT 91.018 79.929 91.064 95.489 ;
        RECT 80.018 90.929 95.552 91.001 ;
        RECT 90.972 79.975 91.018 95.535 ;
        RECT 80.064 90.883 95.598 90.955 ;
        RECT 90.926 80.021 90.972 95.581 ;
        RECT 80.11 90.837 95.644 90.909 ;
        RECT 90.88 80.067 90.926 95.627 ;
        RECT 80.156 90.791 95.69 90.863 ;
        RECT 90.834 80.113 90.88 95.673 ;
        RECT 80.202 90.745 95.736 90.817 ;
        RECT 90.788 80.159 90.834 95.719 ;
        RECT 80.248 90.699 95.782 90.771 ;
        RECT 90.742 80.205 90.788 95.765 ;
        RECT 80.294 90.653 95.828 90.725 ;
        RECT 90.696 80.251 90.742 95.811 ;
        RECT 80.34 90.607 95.874 90.679 ;
        RECT 90.65 80.297 90.696 95.857 ;
        RECT 80.386 90.561 95.92 90.633 ;
        RECT 90.604 80.343 90.65 95.903 ;
        RECT 80.432 90.515 95.966 90.587 ;
        RECT 90.558 80.389 90.604 95.949 ;
        RECT 80.478 90.469 96.012 90.541 ;
        RECT 90.512 80.435 90.558 95.995 ;
        RECT 80.524 90.423 96.058 90.495 ;
        RECT 90.466 80.481 90.512 96.041 ;
        RECT 80.57 90.377 96.104 90.449 ;
        RECT 90.42 80.527 90.466 96.087 ;
        RECT 80.616 90.331 96.15 90.403 ;
        RECT 90.374 80.573 90.42 96.133 ;
        RECT 80.662 90.285 96.196 90.357 ;
        RECT 90.328 80.619 90.374 96.179 ;
        RECT 80.708 90.239 96.242 90.311 ;
        RECT 90.282 80.665 90.328 96.225 ;
        RECT 80.754 90.193 96.288 90.265 ;
        RECT 90.236 80.711 90.282 96.271 ;
        RECT 80.8 90.147 96.334 90.219 ;
        RECT 90.19 80.757 90.236 96.317 ;
        RECT 80.846 90.101 96.38 90.173 ;
        RECT 90.144 80.803 90.19 96.363 ;
        RECT 80.892 90.055 96.426 90.127 ;
        RECT 90.098 80.849 90.144 96.409 ;
        RECT 80.938 90.009 96.472 90.081 ;
        RECT 90.052 80.895 90.098 96.455 ;
        RECT 80.984 89.963 96.518 90.035 ;
        RECT 90.006 80.941 90.052 96.501 ;
        RECT 81.03 89.917 96.564 89.989 ;
        RECT 89.96 80.987 90.006 96.547 ;
        RECT 81.076 89.871 96.61 89.943 ;
        RECT 89.914 81.033 89.96 96.593 ;
        RECT 81.122 89.825 96.656 89.897 ;
        RECT 89.868 81.079 89.914 96.639 ;
        RECT 81.168 89.779 96.702 89.851 ;
        RECT 89.822 81.125 89.868 96.685 ;
        RECT 81.214 89.733 96.748 89.805 ;
        RECT 89.776 81.171 89.822 96.731 ;
        RECT 81.26 89.687 96.794 89.759 ;
        RECT 89.73 81.217 89.776 96.777 ;
        RECT 81.306 89.641 96.84 89.713 ;
        RECT 89.684 81.263 89.73 96.823 ;
        RECT 81.352 89.595 96.886 89.667 ;
        RECT 89.638 81.309 89.684 96.869 ;
        RECT 81.398 89.549 96.932 89.621 ;
        RECT 89.592 81.355 89.638 96.915 ;
        RECT 81.444 89.503 96.978 89.575 ;
        RECT 89.546 81.401 89.592 96.961 ;
        RECT 81.49 89.457 97.03 89.503 ;
        RECT 89.5 81.447 89.546 97.007 ;
        RECT 78.5 92.447 89.5 110 ;
        RECT 81.536 89.411 110 89.5 ;
        RECT 89.494 81.473 89.5 110 ;
        RECT 81.582 89.365 110 89.5 ;
        RECT 89.448 81.499 89.5 110 ;
        RECT 81.628 89.319 110 89.5 ;
        RECT 89.402 81.545 89.5 110 ;
        RECT 81.674 89.273 110 89.5 ;
        RECT 89.356 81.591 89.5 110 ;
        RECT 81.72 89.227 110 89.5 ;
        RECT 89.31 81.637 89.5 110 ;
        RECT 81.766 89.181 110 89.5 ;
        RECT 89.264 81.683 89.5 110 ;
        RECT 81.812 89.135 110 89.5 ;
        RECT 89.218 81.729 89.5 110 ;
        RECT 81.858 89.089 110 89.5 ;
        RECT 89.172 81.775 89.5 110 ;
        RECT 81.904 89.043 110 89.5 ;
        RECT 89.126 81.821 89.5 110 ;
        RECT 81.95 88.997 110 89.5 ;
        RECT 89.08 81.867 89.5 110 ;
        RECT 81.996 88.951 110 89.5 ;
        RECT 89.034 81.913 89.5 110 ;
        RECT 82.042 88.905 110 89.5 ;
        RECT 88.988 81.959 89.5 110 ;
        RECT 82.088 88.859 110 89.5 ;
        RECT 88.942 82.005 89.5 110 ;
        RECT 82.134 88.813 110 89.5 ;
        RECT 88.896 82.051 89.5 110 ;
        RECT 82.18 88.767 110 89.5 ;
        RECT 88.85 82.097 89.5 110 ;
        RECT 82.226 88.721 110 89.5 ;
        RECT 88.804 82.143 89.5 110 ;
        RECT 82.272 88.675 110 89.5 ;
        RECT 88.758 82.189 89.5 110 ;
        RECT 82.318 88.629 110 89.5 ;
        RECT 88.712 82.235 89.5 110 ;
        RECT 82.364 88.583 110 89.5 ;
        RECT 88.666 82.281 89.5 110 ;
        RECT 82.41 88.537 110 89.5 ;
        RECT 88.62 82.327 89.5 110 ;
        RECT 82.456 88.491 110 89.5 ;
        RECT 88.574 82.373 89.5 110 ;
        RECT 82.502 88.445 110 89.5 ;
        RECT 88.528 82.419 89.5 110 ;
        RECT 82.548 88.399 110 89.5 ;
        RECT 88.482 82.465 89.5 110 ;
        RECT 82.594 88.353 110 89.5 ;
        RECT 88.436 82.511 89.5 110 ;
        RECT 82.64 88.307 110 89.5 ;
        RECT 88.39 82.557 89.5 110 ;
        RECT 82.686 88.261 110 89.5 ;
        RECT 88.344 82.603 89.5 110 ;
        RECT 82.732 88.215 110 89.5 ;
        RECT 88.298 82.649 89.5 110 ;
        RECT 82.778 88.169 110 89.5 ;
        RECT 88.252 82.695 89.5 110 ;
        RECT 82.824 88.123 110 89.5 ;
        RECT 88.206 82.741 89.5 110 ;
        RECT 82.87 88.077 110 89.5 ;
        RECT 88.16 82.787 89.5 110 ;
        RECT 82.916 88.031 110 89.5 ;
        RECT 88.114 82.833 89.5 110 ;
        RECT 82.962 87.985 110 89.5 ;
        RECT 88.068 82.879 89.5 110 ;
        RECT 83.008 87.939 110 89.5 ;
        RECT 88.022 82.925 89.5 110 ;
        RECT 83.054 87.893 110 89.5 ;
        RECT 87.976 82.971 89.5 110 ;
        RECT 83.1 87.847 110 89.5 ;
        RECT 87.93 83.017 89.5 110 ;
        RECT 83.146 87.801 110 89.5 ;
        RECT 87.884 83.063 89.5 110 ;
        RECT 83.192 87.755 110 89.5 ;
        RECT 87.838 83.109 89.5 110 ;
        RECT 83.238 87.709 110 89.5 ;
        RECT 87.792 83.155 89.5 110 ;
        RECT 83.284 87.663 110 89.5 ;
        RECT 87.746 83.201 89.5 110 ;
        RECT 83.33 87.617 110 89.5 ;
        RECT 87.7 83.247 89.5 110 ;
        RECT 83.376 87.571 110 89.5 ;
        RECT 87.654 83.293 89.5 110 ;
        RECT 83.422 87.525 110 89.5 ;
        RECT 87.608 83.339 89.5 110 ;
        RECT 83.468 87.479 110 89.5 ;
        RECT 87.562 83.385 89.5 110 ;
        RECT 83.514 87.433 110 89.5 ;
        RECT 87.516 83.431 89.5 110 ;
        RECT 83.56 87.387 110 89.5 ;
        RECT 87.47 83.477 89.5 110 ;
        RECT 83.606 87.341 110 89.5 ;
        RECT 87.424 83.523 89.5 110 ;
        RECT 83.652 87.295 110 89.5 ;
        RECT 87.378 83.569 89.5 110 ;
        RECT 83.698 87.249 110 89.5 ;
        RECT 87.332 83.615 89.5 110 ;
        RECT 83.744 87.203 110 89.5 ;
        RECT 87.286 83.661 89.5 110 ;
        RECT 83.79 87.157 110 89.5 ;
        RECT 87.24 83.707 89.5 110 ;
        RECT 83.836 87.111 110 89.5 ;
        RECT 87.194 83.753 89.5 110 ;
        RECT 83.882 87.065 110 89.5 ;
        RECT 87.148 83.799 89.5 110 ;
        RECT 83.928 87.019 110 89.5 ;
        RECT 87.102 83.845 89.5 110 ;
        RECT 83.974 86.973 110 89.5 ;
        RECT 87.056 83.891 89.5 110 ;
        RECT 84.02 86.927 110 89.5 ;
        RECT 87.01 83.937 89.5 110 ;
        RECT 84.066 86.881 110 89.5 ;
        RECT 86.964 83.983 89.5 110 ;
        RECT 84.112 86.835 110 89.5 ;
        RECT 86.918 84.029 89.5 110 ;
        RECT 84.158 86.789 110 89.5 ;
        RECT 86.872 84.075 89.5 110 ;
        RECT 84.204 86.743 110 89.5 ;
        RECT 86.826 84.121 89.5 110 ;
        RECT 84.25 86.697 110 89.5 ;
        RECT 86.78 84.167 89.5 110 ;
        RECT 84.296 86.651 110 89.5 ;
        RECT 86.734 84.213 89.5 110 ;
        RECT 84.342 86.605 110 89.5 ;
        RECT 86.688 84.259 89.5 110 ;
        RECT 84.388 86.559 110 89.5 ;
        RECT 86.642 84.305 89.5 110 ;
        RECT 84.434 86.513 110 89.5 ;
        RECT 86.596 84.351 89.5 110 ;
        RECT 84.48 86.467 110 89.5 ;
        RECT 86.55 84.397 89.5 110 ;
        RECT 84.526 86.421 110 89.5 ;
        RECT 86.504 84.443 89.5 110 ;
        RECT 84.572 86.375 110 89.5 ;
        RECT 86.458 84.489 89.5 110 ;
        RECT 84.618 86.329 110 89.5 ;
        RECT 86.412 84.535 89.5 110 ;
        RECT 84.664 86.283 110 89.5 ;
        RECT 86.366 84.581 89.5 110 ;
        RECT 84.71 86.237 110 89.5 ;
        RECT 86.32 84.627 89.5 110 ;
        RECT 84.756 86.191 110 89.5 ;
        RECT 86.274 84.673 89.5 110 ;
        RECT 84.802 86.145 110 89.5 ;
        RECT 86.228 84.719 89.5 110 ;
        RECT 84.848 86.099 110 89.5 ;
        RECT 86.182 84.765 89.5 110 ;
        RECT 84.894 86.053 110 89.5 ;
        RECT 86.136 84.811 89.5 110 ;
        RECT 84.94 86.007 110 89.5 ;
        RECT 86.09 84.857 89.5 110 ;
        RECT 84.986 85.961 110 89.5 ;
        RECT 86.044 84.903 89.5 110 ;
        RECT 85.032 85.915 110 89.5 ;
        RECT 85.998 84.949 89.5 110 ;
        RECT 85.078 85.869 110 89.5 ;
        RECT 85.952 84.995 89.5 110 ;
        RECT 85.124 85.823 110 89.5 ;
        RECT 85.906 85.041 89.5 110 ;
        RECT 85.17 85.777 110 89.5 ;
        RECT 85.86 85.087 89.5 110 ;
        RECT 85.216 85.731 110 89.5 ;
        RECT 85.814 85.133 89.5 110 ;
        RECT 85.262 85.685 110 89.5 ;
        RECT 85.768 85.179 89.5 110 ;
        RECT 85.308 85.639 110 89.5 ;
        RECT 85.722 85.225 89.5 110 ;
        RECT 85.354 85.593 110 89.5 ;
        RECT 85.676 85.271 89.5 110 ;
        RECT 85.4 85.547 110 89.5 ;
        RECT 85.63 85.317 89.5 110 ;
        RECT 85.446 85.501 110 89.5 ;
        RECT 85.584 85.363 89.5 110 ;
        RECT 85.492 85.455 110 89.5 ;
        RECT 85.538 85.409 89.5 110 ;
        RECT 10.032 49.46 27 49.508 ;
        RECT 9.986 49.506 26.954 49.554 ;
        RECT 9.94 49.552 26.908 49.6 ;
        RECT 9.894 49.598 26.862 49.646 ;
        RECT 9.848 49.644 26.816 49.692 ;
        RECT 9.802 49.69 26.77 49.738 ;
        RECT 9.756 49.736 26.724 49.784 ;
        RECT 9.71 49.782 26.678 49.83 ;
        RECT 9.664 49.828 26.632 49.876 ;
        RECT 9.618 49.874 26.586 49.922 ;
        RECT 9.572 49.92 26.54 49.968 ;
        RECT 9.526 49.966 26.494 50.014 ;
        RECT 9.48 50.012 26.448 50.06 ;
        RECT 9.434 50.058 26.402 50.106 ;
        RECT 9.388 50.104 26.356 50.152 ;
        RECT 9.342 50.15 26.31 50.198 ;
        RECT 9.296 50.196 26.264 50.244 ;
        RECT 9.25 50.242 26.218 50.29 ;
        RECT 9.204 50.288 26.172 50.336 ;
        RECT 9.158 50.334 26.126 50.382 ;
        RECT 9.112 50.38 26.08 50.428 ;
        RECT 9.066 50.426 26.034 50.474 ;
        RECT 9.02 50.472 25.988 50.52 ;
        RECT 8.974 50.518 25.942 50.566 ;
        RECT 8.928 50.564 25.896 50.612 ;
        RECT 8.882 50.61 25.85 50.658 ;
        RECT 8.836 50.656 25.804 50.704 ;
        RECT 8.79 50.702 25.758 50.75 ;
        RECT 8.744 50.748 25.712 50.796 ;
        RECT 8.698 50.794 25.666 50.842 ;
        RECT 8.652 50.84 25.62 50.888 ;
        RECT 8.606 50.886 25.574 50.934 ;
        RECT 8.56 50.932 25.528 50.98 ;
        RECT 8.514 50.978 25.482 51.026 ;
        RECT 8.468 51.024 25.436 51.072 ;
        RECT 8.422 51.07 25.39 51.118 ;
        RECT 8.376 51.116 25.344 51.164 ;
        RECT 8.33 51.162 25.298 51.21 ;
        RECT 8.284 51.208 25.252 51.256 ;
        RECT 8.238 51.254 25.206 51.302 ;
        RECT 8.192 51.3 25.16 51.348 ;
        RECT 8.146 51.346 25.114 51.394 ;
        RECT 8.1 51.392 25.068 51.44 ;
        RECT 8.054 51.438 25.022 51.486 ;
        RECT 8.008 51.484 24.976 51.532 ;
        RECT 7.962 51.53 24.93 51.578 ;
        RECT 7.916 51.576 24.884 51.624 ;
        RECT 7.87 51.622 24.838 51.67 ;
        RECT 7.824 51.668 24.792 51.716 ;
        RECT 7.778 51.714 24.746 51.762 ;
        RECT 7.732 51.76 24.7 51.808 ;
        RECT 7.686 51.806 24.654 51.854 ;
        RECT 7.64 51.852 24.608 51.9 ;
        RECT 7.594 51.898 24.562 51.946 ;
        RECT 7.548 51.944 24.516 51.992 ;
        RECT 7.502 51.99 24.47 52.038 ;
        RECT 7.456 52.036 24.424 52.084 ;
        RECT 7.41 52.082 24.378 52.13 ;
        RECT 7.364 52.128 24.332 52.176 ;
        RECT 7.318 52.174 24.286 52.222 ;
        RECT 7.272 52.22 24.24 52.268 ;
        RECT 7.226 52.266 24.194 52.314 ;
        RECT 7.18 52.312 24.148 52.36 ;
        RECT 7.134 52.358 24.102 52.406 ;
        RECT 7.088 52.404 24.056 52.452 ;
        RECT 7.042 52.45 24.01 52.498 ;
        RECT 6.996 52.496 23.964 52.544 ;
        RECT 6.95 52.542 23.918 52.59 ;
        RECT 6.904 52.588 23.872 52.636 ;
        RECT 6.858 52.634 23.826 52.682 ;
        RECT 6.812 52.68 23.78 52.728 ;
        RECT 6.766 52.726 23.734 52.774 ;
        RECT 6.72 52.772 23.688 52.82 ;
        RECT 6.674 52.818 23.642 52.866 ;
        RECT 6.628 52.864 23.596 52.912 ;
        RECT 6.582 52.91 23.55 52.958 ;
        RECT 6.536 52.956 23.504 53.004 ;
        RECT 6.49 53.002 23.458 53.05 ;
        RECT 6.444 53.048 23.412 53.096 ;
        RECT 6.398 53.094 23.366 53.142 ;
        RECT 6.352 53.14 23.32 53.188 ;
        RECT 6.306 53.186 23.274 53.234 ;
        RECT 6.26 53.232 23.228 53.28 ;
        RECT 6.214 53.278 23.182 53.326 ;
        RECT 6.168 53.324 23.136 53.372 ;
        RECT 6.122 53.37 23.09 53.418 ;
        RECT 6.076 53.416 23.044 53.464 ;
        RECT 6.03 53.462 22.998 53.51 ;
        RECT 5.984 53.508 22.952 53.556 ;
        RECT 5.938 53.554 22.906 53.602 ;
        RECT 5.892 53.6 22.86 53.648 ;
        RECT 5.846 53.646 22.814 53.694 ;
        RECT 5.8 53.692 22.768 53.74 ;
        RECT 5.754 53.738 22.722 53.786 ;
        RECT 5.708 53.784 22.676 53.832 ;
        RECT 5.662 53.83 22.63 53.878 ;
        RECT 5.616 53.876 22.584 53.924 ;
        RECT 5.57 53.922 22.538 53.97 ;
        RECT 5.524 53.968 22.492 54.016 ;
        RECT 5.478 54.014 22.446 54.062 ;
        RECT 5.432 54.06 22.4 54.108 ;
        RECT 5.386 54.106 22.354 54.154 ;
        RECT 5.34 54.152 22.308 54.2 ;
        RECT 5.294 54.198 22.262 54.246 ;
        RECT 5.248 54.244 22.216 54.292 ;
        RECT 5.202 54.29 22.17 54.338 ;
        RECT 5.156 54.336 22.124 54.384 ;
        RECT 5.11 54.382 22.078 54.43 ;
        RECT 5.064 54.428 22.032 54.476 ;
        RECT 5.018 54.474 21.986 54.522 ;
        RECT 4.972 54.52 21.94 54.568 ;
        RECT 4.926 54.566 21.894 54.614 ;
        RECT 4.88 54.612 21.848 54.66 ;
        RECT 4.834 54.658 21.802 54.706 ;
        RECT 4.788 54.704 21.756 54.752 ;
        RECT 4.742 54.75 21.71 54.798 ;
        RECT 4.696 54.796 21.664 54.844 ;
        RECT 4.65 54.842 21.618 54.89 ;
        RECT 4.604 54.888 21.572 54.936 ;
        RECT 4.558 54.934 21.526 54.982 ;
        RECT 4.512 54.98 21.48 55.028 ;
        RECT 4.466 55.026 21.434 55.074 ;
        RECT 4.42 55.072 21.388 55.12 ;
        RECT 4.374 55.118 21.342 55.166 ;
        RECT 4.328 55.164 21.296 55.212 ;
        RECT 4.282 55.21 21.25 55.258 ;
        RECT 4.236 55.256 21.204 55.304 ;
        RECT 4.19 55.302 21.158 55.35 ;
        RECT 4.144 55.348 21.112 55.396 ;
        RECT 4.098 55.394 21.066 55.442 ;
        RECT 4.052 55.44 21.02 55.488 ;
        RECT 4.006 55.486 20.974 55.534 ;
        RECT 3.96 55.532 20.928 55.58 ;
        RECT 3.914 55.578 20.882 55.626 ;
        RECT 3.868 55.624 20.836 55.672 ;
        RECT 3.822 55.67 20.79 55.718 ;
        RECT 3.776 55.716 20.744 55.764 ;
        RECT 3.73 55.762 20.698 55.81 ;
        RECT 3.684 55.808 20.652 55.856 ;
        RECT 3.638 55.854 20.606 55.902 ;
        RECT 3.592 55.9 20.56 55.948 ;
        RECT 3.546 55.946 20.514 55.994 ;
        RECT 3.5 55.992 20.468 56.04 ;
        RECT 3.5 55.992 20.422 56.086 ;
        RECT 3.5 55.992 20.376 56.132 ;
        RECT 3.5 55.992 20.33 56.178 ;
        RECT 3.5 55.992 20.284 56.224 ;
        RECT 3.5 55.992 20.238 56.27 ;
        RECT 3.5 55.992 20.192 56.316 ;
        RECT 3.5 55.992 20.146 56.362 ;
        RECT 3.5 55.992 20.1 56.408 ;
        RECT 3.5 55.992 20.054 56.454 ;
        RECT 3.5 55.992 20.008 56.5 ;
        RECT 3.5 55.992 19.962 56.546 ;
        RECT 3.5 55.992 19.916 56.592 ;
        RECT 3.5 55.992 19.87 56.638 ;
        RECT 3.5 55.992 19.824 56.684 ;
        RECT 3.5 55.992 19.778 56.73 ;
        RECT 3.5 55.992 19.732 56.776 ;
        RECT 3.5 55.992 19.686 56.822 ;
        RECT 3.5 55.992 19.64 56.868 ;
        RECT 3.5 55.992 19.594 56.914 ;
        RECT 3.5 55.992 19.548 56.96 ;
        RECT 3.5 55.992 19.502 57.006 ;
        RECT 3.5 55.992 19.456 57.052 ;
        RECT 3.5 55.992 19.41 57.098 ;
        RECT 3.5 55.992 19.364 57.144 ;
        RECT 3.5 55.992 19.318 57.19 ;
        RECT 3.5 55.992 19.272 57.236 ;
        RECT 3.5 55.992 19.226 57.282 ;
        RECT 3.5 55.992 19.18 57.328 ;
        RECT 3.5 55.992 19.134 57.374 ;
        RECT 3.5 55.992 19.088 57.42 ;
        RECT 3.5 55.992 19.042 57.466 ;
        RECT 3.5 55.992 18.996 57.512 ;
        RECT 3.5 55.992 18.95 57.558 ;
        RECT 3.5 55.992 18.904 57.604 ;
        RECT 3.5 55.992 18.858 57.65 ;
        RECT 3.5 55.992 18.812 57.696 ;
        RECT 3.5 55.992 18.766 57.742 ;
        RECT 3.5 55.992 18.72 57.788 ;
        RECT 3.5 55.992 18.674 57.834 ;
        RECT 3.5 55.992 18.628 57.88 ;
        RECT 3.5 55.992 18.582 57.926 ;
        RECT 3.5 55.992 18.536 57.972 ;
        RECT 3.5 55.992 18.49 58.018 ;
        RECT 3.5 55.992 18.444 58.064 ;
        RECT 3.5 55.992 18.398 58.11 ;
        RECT 3.5 55.992 18.352 58.156 ;
        RECT 3.5 55.992 18.306 58.202 ;
        RECT 3.5 55.992 18.26 58.248 ;
        RECT 3.5 55.992 18.214 58.294 ;
        RECT 3.5 55.992 18.168 58.34 ;
        RECT 3.5 55.992 18.122 58.386 ;
        RECT 3.5 55.992 18.076 58.432 ;
        RECT 3.5 55.992 18.03 58.478 ;
        RECT 3.5 55.992 17.984 58.524 ;
        RECT 3.5 55.992 17.938 58.57 ;
        RECT 3.5 55.992 17.892 58.616 ;
        RECT 3.5 55.992 17.846 58.662 ;
        RECT 3.5 55.992 17.8 58.708 ;
        RECT 3.5 55.992 17.754 58.754 ;
        RECT 3.5 55.992 17.708 58.8 ;
        RECT 3.5 55.992 17.662 58.846 ;
        RECT 3.5 55.992 17.616 58.892 ;
        RECT 3.5 55.992 17.57 58.938 ;
        RECT 3.5 55.992 17.524 58.984 ;
        RECT 3.5 55.992 17.478 59.03 ;
        RECT 3.5 55.992 17.432 59.076 ;
        RECT 3.5 55.992 17.386 59.122 ;
        RECT 3.5 55.992 17.34 59.168 ;
        RECT 3.5 55.992 17.294 59.214 ;
        RECT 3.5 55.992 17.248 59.26 ;
        RECT 3.5 55.992 17.202 59.306 ;
        RECT 3.5 55.992 17.156 59.352 ;
        RECT 3.5 55.992 17.11 59.398 ;
        RECT 3.5 55.992 17.064 59.444 ;
        RECT 3.5 55.992 17.018 59.49 ;
        RECT 3.5 55.992 16.972 59.536 ;
        RECT 3.5 55.992 16.926 59.582 ;
        RECT 3.5 55.992 16.88 59.628 ;
        RECT 3.5 55.992 16.834 59.674 ;
        RECT 3.5 55.992 16.788 59.72 ;
        RECT 3.5 55.992 16.742 59.766 ;
        RECT 3.5 55.992 16.696 59.812 ;
        RECT 3.5 55.992 16.65 59.858 ;
        RECT 3.5 55.992 16.604 59.904 ;
        RECT 3.5 55.992 16.558 59.95 ;
        RECT 3.5 55.992 16.512 59.996 ;
        RECT 3.5 55.992 16.466 60.042 ;
        RECT 3.5 55.992 16.42 60.088 ;
        RECT 3.5 55.992 16.374 60.134 ;
        RECT 3.5 55.992 16.328 60.18 ;
        RECT 3.5 55.992 16.282 60.226 ;
        RECT 3.5 55.992 16.236 60.272 ;
        RECT 3.5 55.992 16.19 60.318 ;
        RECT 3.5 55.992 16.144 60.364 ;
        RECT 3.5 55.992 16.098 60.41 ;
        RECT 3.5 55.992 16.052 60.456 ;
        RECT 3.5 55.992 16.006 60.502 ;
        RECT 3.5 55.992 15.96 60.548 ;
        RECT 3.5 55.992 15.914 60.594 ;
        RECT 3.5 55.992 15.868 60.64 ;
        RECT 3.5 55.992 15.822 60.686 ;
        RECT 3.5 55.992 15.776 60.732 ;
        RECT 3.5 55.992 15.73 60.778 ;
        RECT 3.5 55.992 15.684 60.824 ;
        RECT 3.5 55.992 15.638 60.87 ;
        RECT 3.5 55.992 15.592 60.916 ;
        RECT 3.5 55.992 15.546 60.962 ;
        RECT 3.5 55.992 15.5 110 ;
        RECT 62.764 17 110 29 ;
        RECT 50.758 28.984 67.733 29.024 ;
        RECT 45.836 33.906 62.765 33.971 ;
        RECT 62.718 17.024 62.764 33.994 ;
        RECT 45.79 33.952 62.718 34.04 ;
        RECT 45.882 33.86 62.811 33.947 ;
        RECT 62.672 17.07 62.718 34.04 ;
        RECT 45.744 33.998 62.672 34.086 ;
        RECT 45.928 33.814 62.857 33.901 ;
        RECT 62.626 17.116 62.672 34.086 ;
        RECT 45.698 34.044 62.626 34.132 ;
        RECT 45.974 33.768 62.903 33.855 ;
        RECT 62.58 17.162 62.626 34.132 ;
        RECT 45.652 34.09 62.58 34.178 ;
        RECT 46.02 33.722 62.949 33.809 ;
        RECT 62.534 17.208 62.58 34.178 ;
        RECT 45.606 34.136 62.534 34.224 ;
        RECT 46.066 33.676 62.995 33.763 ;
        RECT 62.488 17.254 62.534 34.224 ;
        RECT 45.56 34.182 62.488 34.27 ;
        RECT 46.112 33.63 63.041 33.717 ;
        RECT 62.442 17.3 62.488 34.27 ;
        RECT 45.514 34.228 62.442 34.316 ;
        RECT 46.158 33.584 63.087 33.671 ;
        RECT 62.396 17.346 62.442 34.316 ;
        RECT 45.468 34.274 62.396 34.362 ;
        RECT 46.204 33.538 63.133 33.625 ;
        RECT 62.35 17.392 62.396 34.362 ;
        RECT 45.422 34.32 62.35 34.408 ;
        RECT 46.25 33.492 63.179 33.579 ;
        RECT 62.304 17.438 62.35 34.408 ;
        RECT 45.376 34.366 62.304 34.454 ;
        RECT 46.296 33.446 63.225 33.533 ;
        RECT 62.258 17.484 62.304 34.454 ;
        RECT 45.33 34.412 62.258 34.5 ;
        RECT 46.342 33.4 63.271 33.487 ;
        RECT 62.212 17.53 62.258 34.5 ;
        RECT 45.284 34.458 62.212 34.546 ;
        RECT 46.388 33.354 63.317 33.441 ;
        RECT 62.166 17.576 62.212 34.546 ;
        RECT 45.238 34.504 62.166 34.592 ;
        RECT 46.434 33.308 63.363 33.395 ;
        RECT 62.12 17.622 62.166 34.592 ;
        RECT 45.192 34.55 62.12 34.638 ;
        RECT 46.48 33.262 63.409 33.349 ;
        RECT 62.074 17.668 62.12 34.638 ;
        RECT 45.146 34.596 62.074 34.684 ;
        RECT 46.526 33.216 63.455 33.303 ;
        RECT 62.028 17.714 62.074 34.684 ;
        RECT 45.1 34.642 62.028 34.73 ;
        RECT 46.572 33.17 63.501 33.257 ;
        RECT 61.982 17.76 62.028 34.73 ;
        RECT 45.054 34.688 61.982 34.776 ;
        RECT 46.618 33.124 63.547 33.211 ;
        RECT 61.936 17.806 61.982 34.776 ;
        RECT 45.008 34.734 61.936 34.822 ;
        RECT 46.664 33.078 63.593 33.165 ;
        RECT 61.89 17.852 61.936 34.822 ;
        RECT 44.962 34.78 61.89 34.868 ;
        RECT 46.71 33.032 63.639 33.119 ;
        RECT 61.844 17.898 61.89 34.868 ;
        RECT 44.916 34.826 61.844 34.914 ;
        RECT 46.756 32.986 63.685 33.073 ;
        RECT 61.798 17.944 61.844 34.914 ;
        RECT 44.87 34.872 61.798 34.96 ;
        RECT 46.802 32.94 63.731 33.027 ;
        RECT 61.752 17.99 61.798 34.96 ;
        RECT 44.824 34.918 61.752 35.006 ;
        RECT 46.848 32.894 63.777 32.981 ;
        RECT 61.706 18.036 61.752 35.006 ;
        RECT 44.778 34.964 61.706 35.052 ;
        RECT 46.894 32.848 63.823 32.935 ;
        RECT 61.66 18.082 61.706 35.052 ;
        RECT 44.732 35.01 61.66 35.098 ;
        RECT 46.94 32.802 63.869 32.889 ;
        RECT 61.614 18.128 61.66 35.098 ;
        RECT 44.686 35.056 61.614 35.144 ;
        RECT 46.986 32.756 63.915 32.843 ;
        RECT 61.568 18.174 61.614 35.144 ;
        RECT 44.64 35.102 61.568 35.19 ;
        RECT 47.032 32.71 63.961 32.797 ;
        RECT 61.522 18.22 61.568 35.19 ;
        RECT 44.594 35.148 61.522 35.236 ;
        RECT 47.078 32.664 64.007 32.751 ;
        RECT 61.476 18.266 61.522 35.236 ;
        RECT 44.548 35.194 61.476 35.282 ;
        RECT 47.124 32.618 64.053 32.705 ;
        RECT 61.43 18.312 61.476 35.282 ;
        RECT 44.502 35.24 61.43 35.328 ;
        RECT 47.17 32.572 64.099 32.659 ;
        RECT 61.384 18.358 61.43 35.328 ;
        RECT 44.456 35.286 61.384 35.374 ;
        RECT 47.216 32.526 64.145 32.613 ;
        RECT 61.338 18.404 61.384 35.374 ;
        RECT 44.41 35.332 61.338 35.42 ;
        RECT 47.262 32.48 64.191 32.567 ;
        RECT 61.292 18.45 61.338 35.42 ;
        RECT 44.364 35.378 61.292 35.466 ;
        RECT 47.308 32.434 64.237 32.521 ;
        RECT 61.246 18.496 61.292 35.466 ;
        RECT 44.318 35.424 61.246 35.512 ;
        RECT 47.354 32.388 64.283 32.475 ;
        RECT 61.2 18.542 61.246 35.512 ;
        RECT 44.272 35.47 61.2 35.558 ;
        RECT 47.4 32.342 64.329 32.429 ;
        RECT 61.154 18.588 61.2 35.558 ;
        RECT 44.226 35.516 61.154 35.604 ;
        RECT 47.446 32.296 64.375 32.383 ;
        RECT 61.108 18.634 61.154 35.604 ;
        RECT 44.18 35.562 61.108 35.65 ;
        RECT 47.492 32.25 64.421 32.337 ;
        RECT 61.062 18.68 61.108 35.65 ;
        RECT 44.134 35.608 61.062 35.696 ;
        RECT 47.538 32.204 64.467 32.291 ;
        RECT 61.016 18.726 61.062 35.696 ;
        RECT 44.088 35.654 61.016 35.742 ;
        RECT 47.584 32.158 64.513 32.245 ;
        RECT 60.97 18.772 61.016 35.742 ;
        RECT 44.042 35.7 60.97 35.788 ;
        RECT 47.63 32.112 64.559 32.199 ;
        RECT 60.924 18.818 60.97 35.788 ;
        RECT 43.996 35.746 60.924 35.834 ;
        RECT 47.676 32.066 64.605 32.153 ;
        RECT 60.878 18.864 60.924 35.834 ;
        RECT 43.95 35.792 60.878 35.88 ;
        RECT 47.722 32.02 64.651 32.107 ;
        RECT 60.832 18.91 60.878 35.88 ;
        RECT 43.904 35.838 60.832 35.926 ;
        RECT 47.768 31.974 64.697 32.061 ;
        RECT 60.786 18.956 60.832 35.926 ;
        RECT 43.858 35.884 60.786 35.972 ;
        RECT 47.814 31.928 64.743 32.015 ;
        RECT 60.74 19.002 60.786 35.972 ;
        RECT 43.812 35.93 60.74 36.018 ;
        RECT 47.86 31.882 64.789 31.969 ;
        RECT 60.694 19.048 60.74 36.018 ;
        RECT 43.766 35.976 60.694 36.064 ;
        RECT 47.906 31.836 64.835 31.923 ;
        RECT 60.648 19.094 60.694 36.064 ;
        RECT 43.72 36.022 60.648 36.11 ;
        RECT 47.952 31.79 64.881 31.877 ;
        RECT 60.602 19.14 60.648 36.11 ;
        RECT 43.674 36.068 60.602 36.156 ;
        RECT 47.998 31.744 64.927 31.831 ;
        RECT 60.556 19.186 60.602 36.156 ;
        RECT 43.628 36.114 60.556 36.202 ;
        RECT 48.044 31.698 64.973 31.785 ;
        RECT 60.51 19.232 60.556 36.202 ;
        RECT 43.582 36.16 60.51 36.248 ;
        RECT 48.09 31.652 65.019 31.739 ;
        RECT 60.464 19.278 60.51 36.248 ;
        RECT 43.536 36.206 60.464 36.294 ;
        RECT 48.136 31.606 65.065 31.693 ;
        RECT 60.418 19.324 60.464 36.294 ;
        RECT 43.49 36.252 60.418 36.34 ;
        RECT 48.182 31.56 65.111 31.647 ;
        RECT 60.372 19.37 60.418 36.34 ;
        RECT 43.444 36.298 60.372 36.386 ;
        RECT 48.228 31.514 65.157 31.601 ;
        RECT 60.326 19.416 60.372 36.386 ;
        RECT 43.398 36.344 60.326 36.432 ;
        RECT 48.274 31.468 65.203 31.555 ;
        RECT 60.28 19.462 60.326 36.432 ;
        RECT 43.352 36.39 60.28 36.478 ;
        RECT 48.32 31.422 65.249 31.509 ;
        RECT 60.234 19.508 60.28 36.478 ;
        RECT 43.306 36.436 60.234 36.524 ;
        RECT 48.366 31.376 65.295 31.463 ;
        RECT 60.188 19.554 60.234 36.524 ;
        RECT 43.26 36.482 60.188 36.57 ;
        RECT 48.412 31.33 65.341 31.417 ;
        RECT 60.142 19.6 60.188 36.57 ;
        RECT 43.214 36.528 60.142 36.616 ;
        RECT 48.458 31.284 65.387 31.371 ;
        RECT 60.096 19.646 60.142 36.616 ;
        RECT 43.168 36.574 60.096 36.662 ;
        RECT 48.504 31.238 65.433 31.325 ;
        RECT 60.05 19.692 60.096 36.662 ;
        RECT 43.122 36.62 60.05 36.708 ;
        RECT 48.55 31.192 65.479 31.279 ;
        RECT 60.004 19.738 60.05 36.708 ;
        RECT 43.076 36.666 60.004 36.754 ;
        RECT 48.596 31.146 65.525 31.233 ;
        RECT 59.958 19.784 60.004 36.754 ;
        RECT 43.03 36.712 59.958 36.8 ;
        RECT 48.642 31.1 65.571 31.187 ;
        RECT 59.912 19.83 59.958 36.8 ;
        RECT 42.984 36.758 59.912 36.846 ;
        RECT 48.688 31.054 65.617 31.141 ;
        RECT 59.866 19.876 59.912 36.846 ;
        RECT 42.938 36.804 59.866 36.892 ;
        RECT 48.734 31.008 65.663 31.095 ;
        RECT 59.82 19.922 59.866 36.892 ;
        RECT 42.892 36.85 59.82 36.938 ;
        RECT 48.78 30.962 65.709 31.049 ;
        RECT 59.774 19.968 59.82 36.938 ;
        RECT 42.846 36.896 59.774 36.984 ;
        RECT 48.826 30.916 65.755 31.003 ;
        RECT 59.728 20.014 59.774 36.984 ;
        RECT 42.8 36.942 59.728 37.03 ;
        RECT 48.872 30.87 65.801 30.957 ;
        RECT 59.682 20.06 59.728 37.03 ;
        RECT 42.754 36.988 59.682 37.076 ;
        RECT 48.918 30.824 65.847 30.911 ;
        RECT 59.636 20.106 59.682 37.076 ;
        RECT 42.708 37.034 59.636 37.122 ;
        RECT 48.964 30.778 65.893 30.865 ;
        RECT 59.59 20.152 59.636 37.122 ;
        RECT 42.662 37.08 59.59 37.168 ;
        RECT 49.01 30.732 65.939 30.819 ;
        RECT 59.544 20.198 59.59 37.168 ;
        RECT 42.616 37.126 59.544 37.214 ;
        RECT 49.056 30.686 65.985 30.773 ;
        RECT 59.498 20.244 59.544 37.214 ;
        RECT 42.57 37.172 59.498 37.26 ;
        RECT 49.102 30.64 66.031 30.727 ;
        RECT 59.452 20.29 59.498 37.26 ;
        RECT 42.524 37.218 59.452 37.306 ;
        RECT 49.148 30.594 66.077 30.681 ;
        RECT 59.406 20.336 59.452 37.306 ;
        RECT 42.478 37.264 59.406 37.352 ;
        RECT 49.194 30.548 66.123 30.635 ;
        RECT 59.36 20.382 59.406 37.352 ;
        RECT 42.432 37.31 59.36 37.398 ;
        RECT 49.24 30.502 66.169 30.589 ;
        RECT 59.314 20.428 59.36 37.398 ;
        RECT 42.386 37.356 59.314 37.444 ;
        RECT 49.286 30.456 66.215 30.543 ;
        RECT 59.268 20.474 59.314 37.444 ;
        RECT 42.34 37.402 59.268 37.49 ;
        RECT 49.332 30.41 66.261 30.497 ;
        RECT 59.222 20.52 59.268 37.49 ;
        RECT 42.294 37.448 59.222 37.536 ;
        RECT 49.378 30.364 66.307 30.451 ;
        RECT 59.176 20.566 59.222 37.536 ;
        RECT 42.248 37.494 59.176 37.582 ;
        RECT 49.424 30.318 66.353 30.405 ;
        RECT 59.13 20.612 59.176 37.582 ;
        RECT 42.202 37.54 59.13 37.628 ;
        RECT 49.47 30.272 66.399 30.359 ;
        RECT 59.084 20.658 59.13 37.628 ;
        RECT 42.156 37.586 59.084 37.674 ;
        RECT 49.516 30.226 66.445 30.313 ;
        RECT 59.038 20.704 59.084 37.674 ;
        RECT 42.11 37.632 59.038 37.72 ;
        RECT 49.562 30.18 66.491 30.267 ;
        RECT 58.992 20.75 59.038 37.72 ;
        RECT 42.064 37.678 58.992 37.766 ;
        RECT 49.608 30.134 66.537 30.221 ;
        RECT 58.946 20.796 58.992 37.766 ;
        RECT 42.018 37.724 58.946 37.812 ;
        RECT 49.654 30.088 66.583 30.175 ;
        RECT 58.9 20.842 58.946 37.812 ;
        RECT 41.972 37.77 58.9 37.858 ;
        RECT 49.7 30.042 66.629 30.129 ;
        RECT 58.854 20.888 58.9 37.858 ;
        RECT 41.926 37.816 58.854 37.904 ;
        RECT 49.746 29.996 66.675 30.083 ;
        RECT 58.808 20.934 58.854 37.904 ;
        RECT 41.88 37.862 58.808 37.95 ;
        RECT 49.792 29.95 66.721 30.037 ;
        RECT 58.762 20.98 58.808 37.95 ;
        RECT 41.834 37.908 58.762 37.996 ;
        RECT 49.838 29.904 66.767 29.991 ;
        RECT 58.716 21.026 58.762 37.996 ;
        RECT 41.788 37.954 58.716 38.042 ;
        RECT 49.884 29.858 66.813 29.945 ;
        RECT 58.67 21.072 58.716 38.042 ;
        RECT 41.742 38 58.67 38.088 ;
        RECT 49.93 29.812 66.859 29.899 ;
        RECT 58.624 21.118 58.67 38.088 ;
        RECT 41.696 38.046 58.624 38.134 ;
        RECT 49.976 29.766 66.905 29.853 ;
        RECT 58.578 21.164 58.624 38.134 ;
        RECT 41.65 38.092 58.578 38.18 ;
        RECT 50.022 29.72 66.951 29.807 ;
        RECT 58.532 21.21 58.578 38.18 ;
        RECT 41.604 38.138 58.532 38.226 ;
        RECT 50.068 29.674 66.997 29.761 ;
        RECT 58.486 21.256 58.532 38.226 ;
        RECT 41.558 38.184 58.486 38.272 ;
        RECT 50.114 29.628 67.043 29.715 ;
        RECT 58.44 21.302 58.486 38.272 ;
        RECT 41.512 38.23 58.44 38.318 ;
        RECT 50.16 29.582 67.089 29.669 ;
        RECT 58.394 21.348 58.44 38.318 ;
        RECT 41.466 38.276 58.394 38.364 ;
        RECT 50.206 29.536 67.135 29.623 ;
        RECT 58.348 21.394 58.394 38.364 ;
        RECT 41.42 38.322 58.348 38.41 ;
        RECT 50.252 29.49 67.181 29.577 ;
        RECT 58.302 21.44 58.348 38.41 ;
        RECT 41.374 38.368 58.302 38.456 ;
        RECT 50.298 29.444 67.227 29.531 ;
        RECT 58.256 21.486 58.302 38.456 ;
        RECT 41.328 38.414 58.256 38.502 ;
        RECT 50.344 29.398 67.273 29.485 ;
        RECT 58.21 21.532 58.256 38.502 ;
        RECT 41.282 38.46 58.21 38.548 ;
        RECT 50.39 29.352 67.319 29.439 ;
        RECT 58.164 21.578 58.21 38.548 ;
        RECT 41.236 38.506 58.164 38.594 ;
        RECT 50.436 29.306 67.365 29.393 ;
        RECT 58.118 21.624 58.164 38.594 ;
        RECT 41.19 38.552 58.118 38.64 ;
        RECT 50.482 29.26 67.411 29.347 ;
        RECT 58.072 21.67 58.118 38.64 ;
        RECT 41.144 38.598 58.072 38.686 ;
        RECT 50.528 29.214 67.457 29.301 ;
        RECT 58.026 21.716 58.072 38.686 ;
        RECT 41.098 38.644 58.026 38.732 ;
        RECT 50.574 29.168 67.503 29.255 ;
        RECT 57.98 21.762 58.026 38.732 ;
        RECT 41.052 38.69 57.98 38.778 ;
        RECT 50.62 29.122 67.549 29.209 ;
        RECT 57.934 21.808 57.98 38.778 ;
        RECT 41.006 38.736 57.934 38.824 ;
        RECT 50.666 29.076 67.595 29.163 ;
        RECT 57.888 21.854 57.934 38.824 ;
        RECT 40.96 38.782 57.888 38.87 ;
        RECT 50.712 29.03 67.641 29.117 ;
        RECT 57.842 21.9 57.888 38.87 ;
        RECT 40.914 38.828 57.842 38.916 ;
        RECT 50.758 28.984 67.687 29.071 ;
        RECT 57.796 21.946 57.842 38.916 ;
        RECT 40.868 38.874 57.796 38.962 ;
        RECT 50.804 28.938 110 29 ;
        RECT 57.75 21.992 57.796 38.962 ;
        RECT 40.822 38.92 57.75 39.008 ;
        RECT 50.85 28.892 110 29 ;
        RECT 57.704 22.038 57.75 39.008 ;
        RECT 40.776 38.966 57.704 39.054 ;
        RECT 50.896 28.846 110 29 ;
        RECT 57.658 22.084 57.704 39.054 ;
        RECT 40.73 39.012 57.658 39.1 ;
        RECT 50.942 28.8 110 29 ;
        RECT 57.612 22.13 57.658 39.1 ;
        RECT 40.684 39.058 57.612 39.146 ;
        RECT 50.988 28.754 110 29 ;
        RECT 57.566 22.176 57.612 39.146 ;
        RECT 40.638 39.104 57.566 39.192 ;
        RECT 51.034 28.708 110 29 ;
        RECT 57.52 22.222 57.566 39.192 ;
        RECT 40.592 39.15 57.52 39.238 ;
        RECT 51.08 28.662 110 29 ;
        RECT 57.474 22.268 57.52 39.238 ;
        RECT 40.546 39.196 57.474 39.284 ;
        RECT 51.126 28.616 110 29 ;
        RECT 57.428 22.314 57.474 39.284 ;
        RECT 40.5 39.242 57.428 39.33 ;
        RECT 51.172 28.57 110 29 ;
        RECT 57.382 22.36 57.428 39.33 ;
        RECT 40.454 39.288 57.382 39.376 ;
        RECT 51.218 28.524 110 29 ;
        RECT 57.336 22.406 57.382 39.376 ;
        RECT 40.408 39.334 57.336 39.422 ;
        RECT 51.264 28.478 110 29 ;
        RECT 57.29 22.452 57.336 39.422 ;
        RECT 40.362 39.38 57.29 39.468 ;
        RECT 51.31 28.432 110 29 ;
        RECT 57.244 22.498 57.29 39.468 ;
        RECT 40.316 39.426 57.244 39.514 ;
        RECT 51.356 28.386 110 29 ;
        RECT 57.198 22.544 57.244 39.514 ;
        RECT 40.27 39.472 57.198 39.56 ;
        RECT 51.402 28.34 110 29 ;
        RECT 57.152 22.59 57.198 39.56 ;
        RECT 40.224 39.518 57.152 39.606 ;
        RECT 51.448 28.294 110 29 ;
        RECT 57.106 22.636 57.152 39.606 ;
        RECT 40.178 39.564 57.106 39.652 ;
        RECT 51.494 28.248 110 29 ;
        RECT 57.06 22.682 57.106 39.652 ;
        RECT 40.132 39.61 57.06 39.698 ;
        RECT 51.54 28.202 110 29 ;
        RECT 57.014 22.728 57.06 39.698 ;
        RECT 40.086 39.656 57.014 39.744 ;
        RECT 51.586 28.156 110 29 ;
        RECT 56.968 22.774 57.014 39.744 ;
        RECT 40.04 39.702 56.968 39.79 ;
        RECT 51.632 28.11 110 29 ;
        RECT 56.922 22.82 56.968 39.79 ;
        RECT 39.994 39.748 56.922 39.836 ;
        RECT 51.678 28.064 110 29 ;
        RECT 56.876 22.866 56.922 39.836 ;
        RECT 39.948 39.794 56.876 39.882 ;
        RECT 51.724 28.018 110 29 ;
        RECT 56.83 22.912 56.876 39.882 ;
        RECT 39.902 39.84 56.83 39.928 ;
        RECT 51.77 27.972 110 29 ;
        RECT 56.784 22.958 56.83 39.928 ;
        RECT 39.856 39.886 56.784 39.974 ;
        RECT 51.816 27.926 110 29 ;
        RECT 56.738 23.004 56.784 39.974 ;
        RECT 39.81 39.932 56.738 40.02 ;
        RECT 51.862 27.88 110 29 ;
        RECT 56.692 23.05 56.738 40.02 ;
        RECT 39.764 39.978 56.692 40.066 ;
        RECT 51.908 27.834 110 29 ;
        RECT 56.646 23.096 56.692 40.066 ;
        RECT 39.718 40.024 56.646 40.112 ;
        RECT 51.954 27.788 110 29 ;
        RECT 56.6 23.142 56.646 40.112 ;
        RECT 39.672 40.07 56.6 40.158 ;
        RECT 52 27.742 110 29 ;
        RECT 56.554 23.188 56.6 40.158 ;
        RECT 39.626 40.116 56.554 40.204 ;
        RECT 52.046 27.696 110 29 ;
        RECT 56.508 23.234 56.554 40.204 ;
        RECT 39.58 40.162 56.508 40.25 ;
        RECT 52.092 27.65 110 29 ;
        RECT 56.462 23.28 56.508 40.25 ;
        RECT 39.534 40.208 56.462 40.296 ;
        RECT 52.138 27.604 110 29 ;
        RECT 56.416 23.326 56.462 40.296 ;
        RECT 39.488 40.254 56.416 40.342 ;
        RECT 52.184 27.558 110 29 ;
        RECT 56.37 23.372 56.416 40.342 ;
        RECT 39.442 40.3 56.37 40.388 ;
        RECT 52.23 27.512 110 29 ;
        RECT 56.324 23.418 56.37 40.388 ;
        RECT 39.396 40.346 56.324 40.434 ;
        RECT 52.276 27.466 110 29 ;
        RECT 56.278 23.464 56.324 40.434 ;
        RECT 39.35 40.392 56.278 40.48 ;
        RECT 52.322 27.42 110 29 ;
        RECT 56.232 23.51 56.278 40.48 ;
        RECT 39.304 40.438 56.232 40.526 ;
        RECT 52.368 27.374 110 29 ;
        RECT 56.186 23.556 56.232 40.526 ;
        RECT 39.258 40.484 56.186 40.572 ;
        RECT 52.414 27.328 110 29 ;
        RECT 56.14 23.602 56.186 40.572 ;
        RECT 39.212 40.53 56.14 40.618 ;
        RECT 52.46 27.282 110 29 ;
        RECT 56.094 23.648 56.14 40.618 ;
        RECT 39.166 40.576 56.094 40.664 ;
        RECT 52.506 27.236 110 29 ;
        RECT 56.048 23.694 56.094 40.664 ;
        RECT 39.12 40.622 56.048 40.71 ;
        RECT 52.552 27.19 110 29 ;
        RECT 56.002 23.74 56.048 40.71 ;
        RECT 39.074 40.668 56.002 40.756 ;
        RECT 52.598 27.144 110 29 ;
        RECT 55.956 23.786 56.002 40.756 ;
        RECT 39.028 40.714 55.956 40.802 ;
        RECT 52.644 27.098 110 29 ;
        RECT 55.91 23.832 55.956 40.802 ;
        RECT 38.982 40.76 55.91 40.848 ;
        RECT 52.69 27.052 110 29 ;
        RECT 55.864 23.878 55.91 40.848 ;
        RECT 38.936 40.806 55.864 40.894 ;
        RECT 52.736 27.006 110 29 ;
        RECT 55.818 23.924 55.864 40.894 ;
        RECT 38.89 40.852 55.818 40.94 ;
        RECT 52.782 26.96 110 29 ;
        RECT 55.772 23.97 55.818 40.94 ;
        RECT 38.844 40.898 55.772 40.986 ;
        RECT 52.828 26.914 110 29 ;
        RECT 55.726 24.016 55.772 40.986 ;
        RECT 38.798 40.944 55.726 41.032 ;
        RECT 52.874 26.868 110 29 ;
        RECT 55.68 24.062 55.726 41.032 ;
        RECT 38.752 40.99 55.68 41.078 ;
        RECT 52.92 26.822 110 29 ;
        RECT 55.634 24.108 55.68 41.078 ;
        RECT 38.706 41.036 55.634 41.124 ;
        RECT 52.966 26.776 110 29 ;
        RECT 55.588 24.154 55.634 41.124 ;
        RECT 38.66 41.082 55.588 41.17 ;
        RECT 53.012 26.73 110 29 ;
        RECT 55.542 24.2 55.588 41.17 ;
        RECT 38.614 41.128 55.542 41.216 ;
        RECT 53.058 26.684 110 29 ;
        RECT 55.496 24.246 55.542 41.216 ;
        RECT 38.568 41.174 55.496 41.262 ;
        RECT 53.104 26.638 110 29 ;
        RECT 55.45 24.292 55.496 41.262 ;
        RECT 38.522 41.22 55.45 41.308 ;
        RECT 53.15 26.592 110 29 ;
        RECT 55.404 24.338 55.45 41.308 ;
        RECT 38.476 41.266 55.404 41.354 ;
        RECT 53.196 26.546 110 29 ;
        RECT 55.358 24.384 55.404 41.354 ;
        RECT 38.43 41.312 55.358 41.4 ;
        RECT 53.242 26.5 110 29 ;
        RECT 55.312 24.43 55.358 41.4 ;
        RECT 38.384 41.358 55.312 41.446 ;
        RECT 53.288 26.454 110 29 ;
        RECT 55.266 24.476 55.312 41.446 ;
        RECT 38.338 41.404 55.266 41.492 ;
        RECT 53.334 26.408 110 29 ;
        RECT 55.22 24.522 55.266 41.492 ;
        RECT 38.292 41.45 55.22 41.538 ;
        RECT 53.38 26.362 110 29 ;
        RECT 55.174 24.568 55.22 41.538 ;
        RECT 38.246 41.496 55.174 41.584 ;
        RECT 53.426 26.316 110 29 ;
        RECT 55.128 24.614 55.174 41.584 ;
        RECT 38.2 41.542 55.128 41.63 ;
        RECT 53.472 26.27 110 29 ;
        RECT 55.082 24.66 55.128 41.63 ;
        RECT 38.154 41.588 55.082 41.676 ;
        RECT 53.518 26.224 110 29 ;
        RECT 55.036 24.706 55.082 41.676 ;
        RECT 38.108 41.634 55.036 41.722 ;
        RECT 53.564 26.178 110 29 ;
        RECT 54.99 24.752 55.036 41.722 ;
        RECT 38.062 41.68 54.99 41.768 ;
        RECT 53.61 26.132 110 29 ;
        RECT 54.944 24.798 54.99 41.768 ;
        RECT 38.016 41.726 54.944 41.814 ;
        RECT 53.656 26.086 110 29 ;
        RECT 54.898 24.844 54.944 41.814 ;
        RECT 37.97 41.772 54.898 41.86 ;
        RECT 53.702 26.04 110 29 ;
        RECT 54.852 24.89 54.898 41.86 ;
        RECT 37.924 41.818 54.852 41.906 ;
        RECT 53.748 25.994 110 29 ;
        RECT 54.806 24.936 54.852 41.906 ;
        RECT 37.878 41.864 54.806 41.952 ;
        RECT 53.794 25.948 110 29 ;
        RECT 54.76 24.982 54.806 41.952 ;
        RECT 37.832 41.91 54.76 41.998 ;
        RECT 53.84 25.902 110 29 ;
        RECT 54.714 25.028 54.76 41.998 ;
        RECT 37.786 41.956 54.714 42.044 ;
        RECT 53.886 25.856 110 29 ;
        RECT 54.668 25.074 54.714 42.044 ;
        RECT 37.74 42.002 54.668 42.09 ;
        RECT 53.932 25.81 110 29 ;
        RECT 54.622 25.12 54.668 42.09 ;
        RECT 37.694 42.048 54.622 42.136 ;
        RECT 53.978 25.764 110 29 ;
        RECT 54.576 25.166 54.622 42.136 ;
        RECT 37.648 42.094 54.576 42.182 ;
        RECT 54.024 25.718 110 29 ;
        RECT 54.53 25.212 54.576 42.182 ;
        RECT 37.602 42.14 54.53 42.228 ;
        RECT 54.07 25.672 110 29 ;
        RECT 54.484 25.258 54.53 42.228 ;
        RECT 37.556 42.186 54.484 42.274 ;
        RECT 54.116 25.626 110 29 ;
        RECT 54.438 25.304 54.484 42.274 ;
        RECT 37.51 42.232 54.438 42.32 ;
        RECT 54.162 25.58 110 29 ;
        RECT 54.392 25.35 54.438 42.32 ;
        RECT 37.464 42.278 54.392 42.366 ;
        RECT 54.208 25.534 110 29 ;
        RECT 54.346 25.396 54.392 42.366 ;
        RECT 37.418 42.324 54.346 42.412 ;
        RECT 54.254 25.488 110 29 ;
        RECT 54.3 25.442 54.346 42.412 ;
        RECT 37.372 42.37 54.3 42.458 ;
        RECT 37.326 42.416 54.254 42.504 ;
        RECT 37.28 42.462 54.208 42.55 ;
        RECT 37.234 42.508 54.162 42.596 ;
        RECT 37.188 42.554 54.116 42.642 ;
        RECT 37.142 42.6 54.07 42.688 ;
        RECT 37.096 42.646 54.024 42.734 ;
        RECT 37.05 42.692 53.978 42.78 ;
        RECT 37.004 42.738 53.932 42.826 ;
        RECT 36.958 42.784 53.886 42.872 ;
        RECT 36.912 42.83 53.84 42.918 ;
        RECT 36.866 42.876 53.794 42.964 ;
        RECT 36.82 42.922 53.748 43.01 ;
        RECT 36.774 42.968 53.702 43.056 ;
        RECT 36.728 43.014 53.656 43.102 ;
        RECT 36.682 43.06 53.61 43.148 ;
        RECT 36.636 43.106 53.564 43.194 ;
        RECT 36.59 43.152 53.518 43.24 ;
        RECT 36.544 43.198 53.472 43.286 ;
        RECT 36.498 43.244 53.426 43.332 ;
        RECT 36.452 43.29 53.38 43.378 ;
        RECT 36.406 43.336 53.334 43.424 ;
        RECT 36.36 43.382 53.288 43.47 ;
        RECT 36.314 43.428 53.242 43.516 ;
        RECT 36.268 43.474 53.196 43.562 ;
        RECT 36.222 43.52 53.15 43.608 ;
        RECT 36.176 43.566 53.104 43.654 ;
        RECT 36.13 43.612 53.058 43.7 ;
        RECT 36.084 43.658 53.012 43.746 ;
        RECT 36.038 43.704 52.966 43.792 ;
        RECT 35.992 43.75 52.92 43.838 ;
        RECT 35.946 43.796 52.874 43.884 ;
        RECT 35.9 43.842 52.828 43.93 ;
        RECT 35.854 43.888 52.782 43.976 ;
        RECT 35.808 43.934 52.736 44.022 ;
        RECT 35.762 43.98 52.69 44.068 ;
        RECT 35.716 44.026 52.644 44.114 ;
        RECT 35.67 44.072 52.598 44.16 ;
        RECT 35.624 44.118 52.552 44.206 ;
        RECT 35.578 44.164 52.506 44.252 ;
        RECT 35.532 44.21 52.46 44.298 ;
        RECT 35.486 44.256 52.414 44.344 ;
        RECT 35.44 44.302 52.368 44.39 ;
        RECT 35.394 44.348 52.322 44.436 ;
        RECT 35.348 44.394 52.276 44.482 ;
        RECT 35.302 44.44 52.23 44.528 ;
        RECT 35.256 44.486 52.184 44.574 ;
        RECT 35.21 44.532 52.138 44.62 ;
        RECT 35.164 44.578 52.092 44.666 ;
        RECT 35.118 44.624 52.046 44.712 ;
        RECT 35.072 44.67 52 44.758 ;
        RECT 35.026 44.716 51.954 44.804 ;
        RECT 34.98 44.762 51.908 44.85 ;
        RECT 34.934 44.808 51.862 44.896 ;
        RECT 34.888 44.854 51.816 44.942 ;
        RECT 34.842 44.9 51.77 44.988 ;
        RECT 34.796 44.946 51.724 45.034 ;
        RECT 34.75 44.992 51.678 45.08 ;
        RECT 34.704 45.038 51.632 45.126 ;
        RECT 34.658 45.084 51.586 45.172 ;
        RECT 34.612 45.13 51.54 45.218 ;
        RECT 34.566 45.176 51.494 45.264 ;
        RECT 34.52 45.222 51.448 45.31 ;
        RECT 34.474 45.268 51.402 45.356 ;
        RECT 34.428 45.314 51.356 45.402 ;
        RECT 34.382 45.36 51.31 45.448 ;
        RECT 34.336 45.406 51.264 45.494 ;
        RECT 34.29 45.452 51.218 45.54 ;
        RECT 34.244 45.498 51.172 45.586 ;
        RECT 34.198 45.544 51.126 45.632 ;
        RECT 34.152 45.59 51.08 45.678 ;
        RECT 34.106 45.636 51.034 45.724 ;
        RECT 34.06 45.682 50.988 45.77 ;
        RECT 34.014 45.728 50.942 45.816 ;
        RECT 33.968 45.774 50.896 45.862 ;
        RECT 33.922 45.82 50.85 45.908 ;
        RECT 33.876 45.866 50.804 45.954 ;
        RECT 33.83 45.912 50.758 46 ;
        RECT 33.784 45.958 50.712 46.046 ;
        RECT 33.738 46.004 50.666 46.092 ;
        RECT 33.692 46.05 50.62 46.138 ;
        RECT 33.646 46.096 50.574 46.184 ;
        RECT 33.6 46.142 50.528 46.23 ;
        RECT 33.554 46.188 50.482 46.276 ;
        RECT 33.508 46.234 50.436 46.322 ;
        RECT 33.462 46.28 50.39 46.368 ;
        RECT 33.416 46.326 50.344 46.414 ;
        RECT 33.37 46.372 50.298 46.46 ;
        RECT 33.324 46.418 50.252 46.506 ;
        RECT 33.278 46.464 50.206 46.552 ;
        RECT 33.232 46.51 50.16 46.598 ;
        RECT 33.186 46.556 50.114 46.644 ;
        RECT 33.14 46.602 50.068 46.69 ;
        RECT 33.094 46.648 50.022 46.736 ;
        RECT 33.048 46.694 49.976 46.782 ;
        RECT 33.002 46.74 49.93 46.828 ;
        RECT 32.956 46.786 49.884 46.874 ;
        RECT 32.91 46.832 49.838 46.92 ;
        RECT 32.864 46.878 49.792 46.966 ;
        RECT 32.818 46.924 49.746 47.012 ;
        RECT 32.772 46.97 49.7 47.058 ;
        RECT 32.726 47.016 49.654 47.104 ;
        RECT 32.68 47.062 49.608 47.15 ;
        RECT 32.634 47.108 49.562 47.196 ;
        RECT 32.588 47.154 49.516 47.242 ;
        RECT 32.542 47.2 49.47 47.288 ;
        RECT 32.496 47.246 49.424 47.334 ;
        RECT 32.45 47.292 49.378 47.38 ;
        RECT 32.404 47.338 49.332 47.426 ;
        RECT 32.358 47.384 49.286 47.472 ;
        RECT 32.312 47.43 49.24 47.518 ;
        RECT 32.266 47.476 49.194 47.564 ;
        RECT 32.22 47.522 49.148 47.61 ;
        RECT 32.174 47.568 49.102 47.656 ;
        RECT 32.128 47.614 49.056 47.702 ;
        RECT 32.082 47.66 49.01 47.748 ;
        RECT 32.036 47.706 48.964 47.794 ;
        RECT 31.99 47.752 48.918 47.84 ;
        RECT 31.944 47.798 48.872 47.886 ;
        RECT 31.898 47.844 48.826 47.932 ;
        RECT 31.852 47.89 48.78 47.978 ;
        RECT 31.806 47.936 48.734 48.024 ;
        RECT 31.76 47.982 48.688 48.07 ;
        RECT 31.714 48.028 48.642 48.116 ;
        RECT 31.668 48.074 48.596 48.162 ;
        RECT 31.622 48.12 48.55 48.208 ;
        RECT 31.576 48.166 48.504 48.254 ;
        RECT 31.53 48.212 48.458 48.3 ;
        RECT 31.484 48.258 48.412 48.346 ;
        RECT 31.438 48.304 48.366 48.392 ;
        RECT 31.392 48.35 48.32 48.438 ;
        RECT 31.346 48.396 48.274 48.484 ;
        RECT 31.3 48.442 48.228 48.53 ;
        RECT 31.254 48.488 48.182 48.576 ;
        RECT 31.208 48.534 48.136 48.622 ;
        RECT 31.162 48.58 48.09 48.668 ;
        RECT 31.116 48.626 48.044 48.714 ;
        RECT 31.07 48.672 47.998 48.76 ;
        RECT 31.024 48.718 47.952 48.806 ;
        RECT 30.978 48.764 47.906 48.852 ;
        RECT 30.932 48.81 47.86 48.898 ;
        RECT 30.886 48.856 47.814 48.944 ;
        RECT 30.84 48.902 47.768 48.99 ;
        RECT 30.794 48.948 47.722 49.036 ;
        RECT 30.748 48.994 47.676 49.082 ;
        RECT 30.702 49.04 47.63 49.128 ;
        RECT 30.656 49.086 47.584 49.174 ;
        RECT 30.61 49.132 47.538 49.22 ;
        RECT 30.564 49.178 47.492 49.266 ;
        RECT 30.518 49.224 47.446 49.312 ;
        RECT 30.472 49.27 47.4 49.358 ;
        RECT 30.426 49.316 47.354 49.404 ;
        RECT 30.38 49.362 47.308 49.45 ;
        RECT 30.334 49.408 47.262 49.496 ;
        RECT 30.288 49.454 47.216 49.542 ;
        RECT 30.242 49.5 47.17 49.588 ;
        RECT 30.196 49.546 47.124 49.634 ;
        RECT 30.15 49.592 47.078 49.68 ;
        RECT 30.104 49.638 47.032 49.726 ;
        RECT 30.058 49.684 46.986 49.772 ;
        RECT 30.012 49.73 46.94 49.818 ;
        RECT 29.966 49.776 46.894 49.864 ;
        RECT 29.92 49.822 46.848 49.91 ;
        RECT 29.874 49.868 46.802 49.956 ;
        RECT 29.828 49.914 46.756 50.002 ;
        RECT 29.782 49.96 46.71 50.048 ;
        RECT 29.736 50.006 46.664 50.094 ;
        RECT 29.69 50.052 46.618 50.14 ;
        RECT 29.644 50.098 46.572 50.186 ;
        RECT 29.598 50.144 46.526 50.232 ;
        RECT 29.552 50.19 46.48 50.278 ;
        RECT 29.506 50.236 46.434 50.324 ;
        RECT 29.46 50.282 46.388 50.37 ;
        RECT 29.414 50.328 46.342 50.416 ;
        RECT 29.368 50.374 46.296 50.462 ;
        RECT 29.322 50.42 46.25 50.508 ;
        RECT 29.276 50.466 46.204 50.554 ;
        RECT 29.23 50.512 46.158 50.6 ;
        RECT 29.184 50.558 46.112 50.646 ;
        RECT 29.138 50.604 46.066 50.692 ;
        RECT 29.092 50.65 46.02 50.738 ;
        RECT 29 50.742 45.974 50.784 ;
        RECT 29.046 50.696 45.974 50.784 ;
        RECT 28.96 50.785 45.928 50.83 ;
        RECT 28.914 50.828 45.882 50.876 ;
        RECT 28.868 50.874 45.836 50.922 ;
        RECT 28.822 50.92 45.79 50.968 ;
        RECT 28.776 50.966 45.744 51.014 ;
        RECT 28.73 51.012 45.698 51.06 ;
        RECT 28.684 51.058 45.652 51.106 ;
        RECT 28.638 51.104 45.606 51.152 ;
        RECT 28.592 51.15 45.56 51.198 ;
        RECT 28.546 51.196 45.514 51.244 ;
        RECT 28.5 51.242 45.468 51.29 ;
        RECT 28.454 51.288 45.422 51.336 ;
        RECT 28.408 51.334 45.376 51.382 ;
        RECT 56.015 3.5 110 15.5 ;
        RECT 39.052 20.44 56.015 20.488 ;
        RECT 39.098 20.394 56.061 20.447 ;
        RECT 55.98 3.517 56.015 20.488 ;
        RECT 39.144 20.348 56.107 20.401 ;
        RECT 55.934 3.558 55.98 20.528 ;
        RECT 39.006 20.486 55.934 20.574 ;
        RECT 39.19 20.302 56.153 20.355 ;
        RECT 55.888 3.604 55.934 20.574 ;
        RECT 38.96 20.532 55.888 20.62 ;
        RECT 39.236 20.256 56.199 20.309 ;
        RECT 55.842 3.65 55.888 20.62 ;
        RECT 38.914 20.578 55.842 20.666 ;
        RECT 39.282 20.21 56.245 20.263 ;
        RECT 55.796 3.696 55.842 20.666 ;
        RECT 38.868 20.624 55.796 20.712 ;
        RECT 39.328 20.164 56.291 20.217 ;
        RECT 55.75 3.742 55.796 20.712 ;
        RECT 38.822 20.67 55.75 20.758 ;
        RECT 39.374 20.118 56.337 20.171 ;
        RECT 55.704 3.788 55.75 20.758 ;
        RECT 38.776 20.716 55.704 20.804 ;
        RECT 39.42 20.072 56.383 20.125 ;
        RECT 55.658 3.834 55.704 20.804 ;
        RECT 38.73 20.762 55.658 20.85 ;
        RECT 39.466 20.026 56.429 20.079 ;
        RECT 55.612 3.88 55.658 20.85 ;
        RECT 38.684 20.808 55.612 20.896 ;
        RECT 39.512 19.98 56.475 20.033 ;
        RECT 55.566 3.926 55.612 20.896 ;
        RECT 38.638 20.854 55.566 20.942 ;
        RECT 39.558 19.934 56.521 19.987 ;
        RECT 55.52 3.972 55.566 20.942 ;
        RECT 38.592 20.9 55.52 20.988 ;
        RECT 39.604 19.888 56.567 19.941 ;
        RECT 55.474 4.018 55.52 20.988 ;
        RECT 38.546 20.946 55.474 21.034 ;
        RECT 39.65 19.842 56.613 19.895 ;
        RECT 55.428 4.064 55.474 21.034 ;
        RECT 38.5 20.992 55.428 21.08 ;
        RECT 39.696 19.796 56.659 19.849 ;
        RECT 55.382 4.11 55.428 21.08 ;
        RECT 38.454 21.038 55.382 21.126 ;
        RECT 39.742 19.75 56.705 19.803 ;
        RECT 55.336 4.156 55.382 21.126 ;
        RECT 38.408 21.084 55.336 21.172 ;
        RECT 39.788 19.704 56.751 19.757 ;
        RECT 55.29 4.202 55.336 21.172 ;
        RECT 38.362 21.13 55.29 21.218 ;
        RECT 39.834 19.658 56.797 19.711 ;
        RECT 55.244 4.248 55.29 21.218 ;
        RECT 38.316 21.176 55.244 21.264 ;
        RECT 39.88 19.612 56.843 19.665 ;
        RECT 55.198 4.294 55.244 21.264 ;
        RECT 38.27 21.222 55.198 21.31 ;
        RECT 39.926 19.566 56.889 19.619 ;
        RECT 55.152 4.34 55.198 21.31 ;
        RECT 38.224 21.268 55.152 21.356 ;
        RECT 39.972 19.52 56.935 19.573 ;
        RECT 55.106 4.386 55.152 21.356 ;
        RECT 38.178 21.314 55.106 21.402 ;
        RECT 40.018 19.474 56.981 19.527 ;
        RECT 55.06 4.432 55.106 21.402 ;
        RECT 38.132 21.36 55.06 21.448 ;
        RECT 40.064 19.428 57.027 19.481 ;
        RECT 55.014 4.478 55.06 21.448 ;
        RECT 38.086 21.406 55.014 21.494 ;
        RECT 40.11 19.382 57.073 19.435 ;
        RECT 54.968 4.524 55.014 21.494 ;
        RECT 38.04 21.452 54.968 21.54 ;
        RECT 40.156 19.336 57.119 19.389 ;
        RECT 54.922 4.57 54.968 21.54 ;
        RECT 37.994 21.498 54.922 21.586 ;
        RECT 40.202 19.29 57.165 19.343 ;
        RECT 54.876 4.616 54.922 21.586 ;
        RECT 37.948 21.544 54.876 21.632 ;
        RECT 40.248 19.244 57.211 19.297 ;
        RECT 54.83 4.662 54.876 21.632 ;
        RECT 37.902 21.59 54.83 21.678 ;
        RECT 40.294 19.198 57.257 19.251 ;
        RECT 54.784 4.708 54.83 21.678 ;
        RECT 37.856 21.636 54.784 21.724 ;
        RECT 40.34 19.152 57.303 19.205 ;
        RECT 54.738 4.754 54.784 21.724 ;
        RECT 37.81 21.682 54.738 21.77 ;
        RECT 40.386 19.106 57.349 19.159 ;
        RECT 54.692 4.8 54.738 21.77 ;
        RECT 37.764 21.728 54.692 21.816 ;
        RECT 40.432 19.06 57.395 19.113 ;
        RECT 54.646 4.846 54.692 21.816 ;
        RECT 37.718 21.774 54.646 21.862 ;
        RECT 40.478 19.014 57.441 19.067 ;
        RECT 54.6 4.892 54.646 21.862 ;
        RECT 37.672 21.82 54.6 21.908 ;
        RECT 40.524 18.968 57.487 19.021 ;
        RECT 54.554 4.938 54.6 21.908 ;
        RECT 37.626 21.866 54.554 21.954 ;
        RECT 40.57 18.922 57.533 18.975 ;
        RECT 54.508 4.984 54.554 21.954 ;
        RECT 37.58 21.912 54.508 22 ;
        RECT 40.616 18.876 57.579 18.929 ;
        RECT 54.462 5.03 54.508 22 ;
        RECT 37.534 21.958 54.462 22.046 ;
        RECT 40.662 18.83 57.625 18.883 ;
        RECT 54.416 5.076 54.462 22.046 ;
        RECT 37.488 22.004 54.416 22.092 ;
        RECT 40.708 18.784 57.671 18.837 ;
        RECT 54.37 5.122 54.416 22.092 ;
        RECT 37.442 22.05 54.37 22.138 ;
        RECT 40.754 18.738 57.717 18.791 ;
        RECT 54.324 5.168 54.37 22.138 ;
        RECT 37.396 22.096 54.324 22.184 ;
        RECT 40.8 18.692 57.763 18.745 ;
        RECT 54.278 5.214 54.324 22.184 ;
        RECT 37.35 22.142 54.278 22.23 ;
        RECT 40.846 18.646 57.809 18.699 ;
        RECT 54.232 5.26 54.278 22.23 ;
        RECT 37.304 22.188 54.232 22.276 ;
        RECT 40.892 18.6 57.855 18.653 ;
        RECT 54.186 5.306 54.232 22.276 ;
        RECT 37.258 22.234 54.186 22.322 ;
        RECT 40.938 18.554 57.901 18.607 ;
        RECT 54.14 5.352 54.186 22.322 ;
        RECT 37.212 22.28 54.14 22.368 ;
        RECT 40.984 18.508 57.947 18.561 ;
        RECT 54.094 5.398 54.14 22.368 ;
        RECT 37.166 22.326 54.094 22.414 ;
        RECT 41.03 18.462 57.993 18.515 ;
        RECT 54.048 5.444 54.094 22.414 ;
        RECT 37.12 22.372 54.048 22.46 ;
        RECT 41.076 18.416 58.039 18.469 ;
        RECT 54.002 5.49 54.048 22.46 ;
        RECT 37.074 22.418 54.002 22.506 ;
        RECT 41.122 18.37 58.085 18.423 ;
        RECT 53.956 5.536 54.002 22.506 ;
        RECT 37.028 22.464 53.956 22.552 ;
        RECT 41.168 18.324 58.131 18.377 ;
        RECT 53.91 5.582 53.956 22.552 ;
        RECT 36.982 22.51 53.91 22.598 ;
        RECT 41.214 18.278 58.177 18.331 ;
        RECT 53.864 5.628 53.91 22.598 ;
        RECT 36.936 22.556 53.864 22.644 ;
        RECT 41.26 18.232 58.223 18.285 ;
        RECT 53.818 5.674 53.864 22.644 ;
        RECT 36.89 22.602 53.818 22.69 ;
        RECT 41.306 18.186 58.269 18.239 ;
        RECT 53.772 5.72 53.818 22.69 ;
        RECT 36.844 22.648 53.772 22.736 ;
        RECT 41.352 18.14 58.315 18.193 ;
        RECT 53.726 5.766 53.772 22.736 ;
        RECT 36.798 22.694 53.726 22.782 ;
        RECT 41.398 18.094 58.361 18.147 ;
        RECT 53.68 5.812 53.726 22.782 ;
        RECT 36.752 22.74 53.68 22.828 ;
        RECT 41.444 18.048 58.407 18.101 ;
        RECT 53.634 5.858 53.68 22.828 ;
        RECT 36.706 22.786 53.634 22.874 ;
        RECT 41.49 18.002 58.453 18.055 ;
        RECT 53.588 5.904 53.634 22.874 ;
        RECT 36.66 22.832 53.588 22.92 ;
        RECT 41.536 17.956 58.499 18.009 ;
        RECT 53.542 5.95 53.588 22.92 ;
        RECT 36.614 22.878 53.542 22.966 ;
        RECT 41.582 17.91 58.545 17.963 ;
        RECT 53.496 5.996 53.542 22.966 ;
        RECT 36.568 22.924 53.496 23.012 ;
        RECT 41.628 17.864 58.591 17.917 ;
        RECT 53.45 6.042 53.496 23.012 ;
        RECT 36.522 22.97 53.45 23.058 ;
        RECT 41.674 17.818 58.637 17.871 ;
        RECT 53.404 6.088 53.45 23.058 ;
        RECT 36.476 23.016 53.404 23.104 ;
        RECT 41.72 17.772 58.683 17.825 ;
        RECT 53.358 6.134 53.404 23.104 ;
        RECT 36.43 23.062 53.358 23.15 ;
        RECT 41.766 17.726 58.729 17.779 ;
        RECT 53.312 6.18 53.358 23.15 ;
        RECT 36.384 23.108 53.312 23.196 ;
        RECT 41.812 17.68 58.775 17.733 ;
        RECT 53.266 6.226 53.312 23.196 ;
        RECT 36.338 23.154 53.266 23.242 ;
        RECT 41.858 17.634 58.821 17.687 ;
        RECT 53.22 6.272 53.266 23.242 ;
        RECT 36.292 23.2 53.22 23.288 ;
        RECT 41.904 17.588 58.867 17.641 ;
        RECT 53.174 6.318 53.22 23.288 ;
        RECT 36.246 23.246 53.174 23.334 ;
        RECT 41.95 17.542 58.913 17.595 ;
        RECT 53.128 6.364 53.174 23.334 ;
        RECT 36.2 23.292 53.128 23.38 ;
        RECT 41.996 17.496 58.959 17.549 ;
        RECT 53.082 6.41 53.128 23.38 ;
        RECT 36.154 23.338 53.082 23.426 ;
        RECT 42.042 17.45 59.005 17.503 ;
        RECT 53.036 6.456 53.082 23.426 ;
        RECT 36.108 23.384 53.036 23.472 ;
        RECT 42.088 17.404 59.051 17.457 ;
        RECT 52.99 6.502 53.036 23.472 ;
        RECT 36.062 23.43 52.99 23.518 ;
        RECT 42.134 17.358 59.097 17.411 ;
        RECT 52.944 6.548 52.99 23.518 ;
        RECT 36.016 23.476 52.944 23.564 ;
        RECT 42.18 17.312 59.143 17.365 ;
        RECT 52.898 6.594 52.944 23.564 ;
        RECT 35.97 23.522 52.898 23.61 ;
        RECT 42.226 17.266 59.189 17.319 ;
        RECT 52.852 6.64 52.898 23.61 ;
        RECT 35.924 23.568 52.852 23.656 ;
        RECT 42.272 17.22 59.235 17.273 ;
        RECT 52.806 6.686 52.852 23.656 ;
        RECT 35.878 23.614 52.806 23.702 ;
        RECT 42.318 17.174 59.281 17.227 ;
        RECT 52.76 6.732 52.806 23.702 ;
        RECT 35.832 23.66 52.76 23.748 ;
        RECT 42.364 17.128 59.327 17.181 ;
        RECT 52.714 6.778 52.76 23.748 ;
        RECT 35.786 23.706 52.714 23.794 ;
        RECT 42.41 17.082 59.373 17.135 ;
        RECT 52.668 6.824 52.714 23.794 ;
        RECT 35.74 23.752 52.668 23.84 ;
        RECT 42.456 17.036 59.419 17.089 ;
        RECT 52.622 6.87 52.668 23.84 ;
        RECT 35.694 23.798 52.622 23.886 ;
        RECT 42.502 16.99 59.465 17.043 ;
        RECT 52.576 6.916 52.622 23.886 ;
        RECT 35.648 23.844 52.576 23.932 ;
        RECT 42.548 16.944 59.511 16.997 ;
        RECT 52.53 6.962 52.576 23.932 ;
        RECT 35.602 23.89 52.53 23.978 ;
        RECT 42.594 16.898 59.557 16.951 ;
        RECT 52.484 7.008 52.53 23.978 ;
        RECT 35.556 23.936 52.484 24.024 ;
        RECT 42.64 16.852 59.603 16.905 ;
        RECT 52.438 7.054 52.484 24.024 ;
        RECT 35.51 23.982 52.438 24.07 ;
        RECT 42.686 16.806 59.649 16.859 ;
        RECT 52.392 7.1 52.438 24.07 ;
        RECT 35.464 24.028 52.392 24.116 ;
        RECT 42.732 16.76 59.695 16.813 ;
        RECT 52.346 7.146 52.392 24.116 ;
        RECT 35.418 24.074 52.346 24.162 ;
        RECT 42.778 16.714 59.741 16.767 ;
        RECT 52.3 7.192 52.346 24.162 ;
        RECT 35.372 24.12 52.3 24.208 ;
        RECT 42.824 16.668 59.787 16.721 ;
        RECT 52.254 7.238 52.3 24.208 ;
        RECT 35.326 24.166 52.254 24.254 ;
        RECT 42.87 16.622 59.833 16.675 ;
        RECT 52.208 7.284 52.254 24.254 ;
        RECT 35.28 24.212 52.208 24.3 ;
        RECT 42.916 16.576 59.879 16.629 ;
        RECT 52.162 7.33 52.208 24.3 ;
        RECT 35.234 24.258 52.162 24.346 ;
        RECT 42.962 16.53 59.925 16.583 ;
        RECT 52.116 7.376 52.162 24.346 ;
        RECT 35.188 24.304 52.116 24.392 ;
        RECT 43.008 16.484 59.971 16.537 ;
        RECT 52.07 7.422 52.116 24.392 ;
        RECT 35.142 24.35 52.07 24.438 ;
        RECT 43.054 16.438 60.017 16.491 ;
        RECT 52.024 7.468 52.07 24.438 ;
        RECT 35.096 24.396 52.024 24.484 ;
        RECT 43.1 16.392 60.063 16.445 ;
        RECT 51.978 7.514 52.024 24.484 ;
        RECT 35.05 24.442 51.978 24.53 ;
        RECT 43.146 16.346 60.109 16.399 ;
        RECT 51.932 7.56 51.978 24.53 ;
        RECT 35.004 24.488 51.932 24.576 ;
        RECT 43.192 16.3 60.155 16.353 ;
        RECT 51.886 7.606 51.932 24.576 ;
        RECT 34.958 24.534 51.886 24.622 ;
        RECT 43.238 16.254 60.201 16.307 ;
        RECT 51.84 7.652 51.886 24.622 ;
        RECT 34.912 24.58 51.84 24.668 ;
        RECT 43.284 16.208 60.247 16.261 ;
        RECT 51.794 7.698 51.84 24.668 ;
        RECT 34.866 24.626 51.794 24.714 ;
        RECT 43.33 16.162 60.293 16.215 ;
        RECT 51.748 7.744 51.794 24.714 ;
        RECT 34.82 24.672 51.748 24.76 ;
        RECT 43.376 16.116 60.339 16.169 ;
        RECT 51.702 7.79 51.748 24.76 ;
        RECT 34.774 24.718 51.702 24.806 ;
        RECT 43.422 16.07 60.385 16.123 ;
        RECT 51.656 7.836 51.702 24.806 ;
        RECT 34.728 24.764 51.656 24.852 ;
        RECT 43.468 16.024 60.431 16.077 ;
        RECT 51.61 7.882 51.656 24.852 ;
        RECT 34.682 24.81 51.61 24.898 ;
        RECT 43.514 15.978 60.477 16.031 ;
        RECT 51.564 7.928 51.61 24.898 ;
        RECT 34.636 24.856 51.564 24.944 ;
        RECT 43.56 15.932 60.523 15.985 ;
        RECT 51.518 7.974 51.564 24.944 ;
        RECT 34.59 24.902 51.518 24.99 ;
        RECT 43.606 15.886 60.569 15.939 ;
        RECT 51.472 8.02 51.518 24.99 ;
        RECT 34.544 24.948 51.472 25.036 ;
        RECT 43.652 15.84 60.615 15.893 ;
        RECT 51.426 8.066 51.472 25.036 ;
        RECT 34.498 24.994 51.426 25.082 ;
        RECT 43.698 15.794 60.661 15.847 ;
        RECT 51.38 8.112 51.426 25.082 ;
        RECT 34.452 25.04 51.38 25.128 ;
        RECT 43.744 15.748 60.707 15.801 ;
        RECT 51.334 8.158 51.38 25.128 ;
        RECT 34.406 25.086 51.334 25.174 ;
        RECT 43.79 15.702 60.753 15.755 ;
        RECT 51.288 8.204 51.334 25.174 ;
        RECT 34.36 25.132 51.288 25.22 ;
        RECT 43.836 15.656 60.799 15.709 ;
        RECT 51.242 8.25 51.288 25.22 ;
        RECT 34.314 25.178 51.242 25.266 ;
        RECT 43.882 15.61 60.845 15.663 ;
        RECT 51.196 8.296 51.242 25.266 ;
        RECT 34.268 25.224 51.196 25.312 ;
        RECT 43.928 15.564 60.891 15.617 ;
        RECT 51.15 8.342 51.196 25.312 ;
        RECT 34.222 25.27 51.15 25.358 ;
        RECT 43.974 15.518 60.937 15.571 ;
        RECT 51.104 8.388 51.15 25.358 ;
        RECT 34.176 25.316 51.104 25.404 ;
        RECT 44.02 15.472 60.983 15.524 ;
        RECT 51.058 8.434 51.104 25.404 ;
        RECT 34.13 25.362 51.058 25.45 ;
        RECT 44.066 15.426 110 15.5 ;
        RECT 51.012 8.48 51.058 25.45 ;
        RECT 34.084 25.408 51.012 25.496 ;
        RECT 44.112 15.38 110 15.5 ;
        RECT 50.966 8.526 51.012 25.496 ;
        RECT 34.038 25.454 50.966 25.542 ;
        RECT 44.158 15.334 110 15.5 ;
        RECT 50.92 8.572 50.966 25.542 ;
        RECT 33.992 25.5 50.92 25.588 ;
        RECT 44.204 15.288 110 15.5 ;
        RECT 50.874 8.618 50.92 25.588 ;
        RECT 33.946 25.546 50.874 25.634 ;
        RECT 44.25 15.242 110 15.5 ;
        RECT 50.828 8.664 50.874 25.634 ;
        RECT 33.9 25.592 50.828 25.68 ;
        RECT 44.296 15.196 110 15.5 ;
        RECT 50.782 8.71 50.828 25.68 ;
        RECT 33.854 25.638 50.782 25.726 ;
        RECT 44.342 15.15 110 15.5 ;
        RECT 50.736 8.756 50.782 25.726 ;
        RECT 33.808 25.684 50.736 25.772 ;
        RECT 44.388 15.104 110 15.5 ;
        RECT 50.69 8.802 50.736 25.772 ;
        RECT 33.762 25.73 50.69 25.818 ;
        RECT 44.434 15.058 110 15.5 ;
        RECT 50.644 8.848 50.69 25.818 ;
        RECT 33.716 25.776 50.644 25.864 ;
        RECT 44.48 15.012 110 15.5 ;
        RECT 50.598 8.894 50.644 25.864 ;
        RECT 33.67 25.822 50.598 25.91 ;
        RECT 44.526 14.966 110 15.5 ;
        RECT 50.552 8.94 50.598 25.91 ;
        RECT 33.624 25.868 50.552 25.956 ;
        RECT 44.572 14.92 110 15.5 ;
        RECT 50.506 8.986 50.552 25.956 ;
        RECT 33.578 25.914 50.506 26.002 ;
        RECT 44.618 14.874 110 15.5 ;
        RECT 50.46 9.032 50.506 26.002 ;
        RECT 33.532 25.96 50.46 26.048 ;
        RECT 44.664 14.828 110 15.5 ;
        RECT 50.414 9.078 50.46 26.048 ;
        RECT 33.486 26.006 50.414 26.094 ;
        RECT 44.71 14.782 110 15.5 ;
        RECT 50.368 9.124 50.414 26.094 ;
        RECT 33.44 26.052 50.368 26.14 ;
        RECT 44.756 14.736 110 15.5 ;
        RECT 50.322 9.17 50.368 26.14 ;
        RECT 33.394 26.098 50.322 26.186 ;
        RECT 44.802 14.69 110 15.5 ;
        RECT 50.276 9.216 50.322 26.186 ;
        RECT 33.348 26.144 50.276 26.232 ;
        RECT 44.848 14.644 110 15.5 ;
        RECT 50.23 9.262 50.276 26.232 ;
        RECT 33.302 26.19 50.23 26.278 ;
        RECT 44.894 14.598 110 15.5 ;
        RECT 50.184 9.308 50.23 26.278 ;
        RECT 33.256 26.236 50.184 26.324 ;
        RECT 44.94 14.552 110 15.5 ;
        RECT 50.138 9.354 50.184 26.324 ;
        RECT 33.21 26.282 50.138 26.37 ;
        RECT 44.986 14.506 110 15.5 ;
        RECT 50.092 9.4 50.138 26.37 ;
        RECT 33.164 26.328 50.092 26.416 ;
        RECT 45.032 14.46 110 15.5 ;
        RECT 50.046 9.446 50.092 26.416 ;
        RECT 33.118 26.374 50.046 26.462 ;
        RECT 45.078 14.414 110 15.5 ;
        RECT 50 9.492 50.046 26.462 ;
        RECT 33.072 26.42 50 26.508 ;
        RECT 45.124 14.368 110 15.5 ;
        RECT 49.954 9.538 50 26.508 ;
        RECT 33.026 26.466 49.954 26.554 ;
        RECT 45.17 14.322 110 15.5 ;
        RECT 49.908 9.584 49.954 26.554 ;
        RECT 32.98 26.512 49.908 26.6 ;
        RECT 45.216 14.276 110 15.5 ;
        RECT 49.862 9.63 49.908 26.6 ;
        RECT 32.934 26.558 49.862 26.646 ;
        RECT 45.262 14.23 110 15.5 ;
        RECT 49.816 9.676 49.862 26.646 ;
        RECT 32.888 26.604 49.816 26.692 ;
        RECT 45.308 14.184 110 15.5 ;
        RECT 49.77 9.722 49.816 26.692 ;
        RECT 32.842 26.65 49.77 26.738 ;
        RECT 45.354 14.138 110 15.5 ;
        RECT 49.724 9.768 49.77 26.738 ;
        RECT 32.796 26.696 49.724 26.784 ;
        RECT 45.4 14.092 110 15.5 ;
        RECT 49.678 9.814 49.724 26.784 ;
        RECT 32.75 26.742 49.678 26.83 ;
        RECT 45.446 14.046 110 15.5 ;
        RECT 49.632 9.86 49.678 26.83 ;
        RECT 32.704 26.788 49.632 26.876 ;
        RECT 45.492 14 110 15.5 ;
        RECT 49.586 9.906 49.632 26.876 ;
        RECT 32.658 26.834 49.586 26.922 ;
        RECT 45.538 13.954 110 15.5 ;
        RECT 49.54 9.952 49.586 26.922 ;
        RECT 32.612 26.88 49.54 26.968 ;
        RECT 45.584 13.908 110 15.5 ;
        RECT 49.494 9.998 49.54 26.968 ;
        RECT 32.566 26.926 49.494 27.014 ;
        RECT 45.63 13.862 110 15.5 ;
        RECT 49.448 10.044 49.494 27.014 ;
        RECT 32.52 26.972 49.448 27.06 ;
        RECT 45.676 13.816 110 15.5 ;
        RECT 49.402 10.09 49.448 27.06 ;
        RECT 32.474 27.018 49.402 27.106 ;
        RECT 45.722 13.77 110 15.5 ;
        RECT 49.356 10.136 49.402 27.106 ;
        RECT 32.428 27.064 49.356 27.152 ;
        RECT 45.768 13.724 110 15.5 ;
        RECT 49.31 10.182 49.356 27.152 ;
        RECT 32.382 27.11 49.31 27.198 ;
        RECT 45.814 13.678 110 15.5 ;
        RECT 49.264 10.228 49.31 27.198 ;
        RECT 32.336 27.156 49.264 27.244 ;
        RECT 45.86 13.632 110 15.5 ;
        RECT 49.218 10.274 49.264 27.244 ;
        RECT 32.29 27.202 49.218 27.29 ;
        RECT 45.906 13.586 110 15.5 ;
        RECT 49.172 10.32 49.218 27.29 ;
        RECT 32.244 27.248 49.172 27.336 ;
        RECT 45.952 13.54 110 15.5 ;
        RECT 49.126 10.366 49.172 27.336 ;
        RECT 32.198 27.294 49.126 27.382 ;
        RECT 45.998 13.494 110 15.5 ;
        RECT 49.08 10.412 49.126 27.382 ;
        RECT 32.152 27.34 49.08 27.428 ;
        RECT 46.044 13.448 110 15.5 ;
        RECT 49.034 10.458 49.08 27.428 ;
        RECT 32.106 27.386 49.034 27.474 ;
        RECT 46.09 13.402 110 15.5 ;
        RECT 48.988 10.504 49.034 27.474 ;
        RECT 32.06 27.432 48.988 27.52 ;
        RECT 46.136 13.356 110 15.5 ;
        RECT 48.942 10.55 48.988 27.52 ;
        RECT 32.014 27.478 48.942 27.566 ;
        RECT 46.182 13.31 110 15.5 ;
        RECT 48.896 10.596 48.942 27.566 ;
        RECT 31.968 27.524 48.896 27.612 ;
        RECT 46.228 13.264 110 15.5 ;
        RECT 48.85 10.642 48.896 27.612 ;
        RECT 31.922 27.57 48.85 27.658 ;
        RECT 46.274 13.218 110 15.5 ;
        RECT 48.804 10.688 48.85 27.658 ;
        RECT 31.876 27.616 48.804 27.704 ;
        RECT 46.32 13.172 110 15.5 ;
        RECT 48.758 10.734 48.804 27.704 ;
        RECT 31.83 27.662 48.758 27.75 ;
        RECT 46.366 13.126 110 15.5 ;
        RECT 48.712 10.78 48.758 27.75 ;
        RECT 31.784 27.708 48.712 27.796 ;
        RECT 46.412 13.08 110 15.5 ;
        RECT 48.666 10.826 48.712 27.796 ;
        RECT 31.738 27.754 48.666 27.842 ;
        RECT 46.458 13.034 110 15.5 ;
        RECT 48.62 10.872 48.666 27.842 ;
        RECT 31.692 27.8 48.62 27.888 ;
        RECT 46.504 12.988 110 15.5 ;
        RECT 48.574 10.918 48.62 27.888 ;
        RECT 31.646 27.846 48.574 27.934 ;
        RECT 46.55 12.942 110 15.5 ;
        RECT 48.528 10.964 48.574 27.934 ;
        RECT 31.6 27.892 48.528 27.98 ;
        RECT 46.596 12.896 110 15.5 ;
        RECT 48.482 11.01 48.528 27.98 ;
        RECT 31.554 27.938 48.482 28.026 ;
        RECT 46.642 12.85 110 15.5 ;
        RECT 48.436 11.056 48.482 28.026 ;
        RECT 31.508 27.984 48.436 28.072 ;
        RECT 46.688 12.804 110 15.5 ;
        RECT 48.39 11.102 48.436 28.072 ;
        RECT 31.462 28.03 48.39 28.118 ;
        RECT 46.734 12.758 110 15.5 ;
        RECT 48.344 11.148 48.39 28.118 ;
        RECT 31.416 28.076 48.344 28.164 ;
        RECT 46.78 12.712 110 15.5 ;
        RECT 48.298 11.194 48.344 28.164 ;
        RECT 31.37 28.122 48.298 28.21 ;
        RECT 46.826 12.666 110 15.5 ;
        RECT 48.252 11.24 48.298 28.21 ;
        RECT 31.324 28.168 48.252 28.256 ;
        RECT 46.872 12.62 110 15.5 ;
        RECT 48.206 11.286 48.252 28.256 ;
        RECT 31.278 28.214 48.206 28.302 ;
        RECT 46.918 12.574 110 15.5 ;
        RECT 48.16 11.332 48.206 28.302 ;
        RECT 31.232 28.26 48.16 28.348 ;
        RECT 46.964 12.528 110 15.5 ;
        RECT 48.114 11.378 48.16 28.348 ;
        RECT 31.186 28.306 48.114 28.394 ;
        RECT 47.01 12.482 110 15.5 ;
        RECT 48.068 11.424 48.114 28.394 ;
        RECT 31.14 28.352 48.068 28.44 ;
        RECT 47.056 12.436 110 15.5 ;
        RECT 48.022 11.47 48.068 28.44 ;
        RECT 31.094 28.398 48.022 28.486 ;
        RECT 47.102 12.39 110 15.5 ;
        RECT 47.976 11.516 48.022 28.486 ;
        RECT 31.048 28.444 47.976 28.532 ;
        RECT 47.148 12.344 110 15.5 ;
        RECT 47.93 11.562 47.976 28.532 ;
        RECT 31.002 28.49 47.93 28.578 ;
        RECT 47.194 12.298 110 15.5 ;
        RECT 47.884 11.608 47.93 28.578 ;
        RECT 30.956 28.536 47.884 28.624 ;
        RECT 47.24 12.252 110 15.5 ;
        RECT 47.838 11.654 47.884 28.624 ;
        RECT 30.91 28.582 47.838 28.67 ;
        RECT 47.286 12.206 110 15.5 ;
        RECT 47.792 11.7 47.838 28.67 ;
        RECT 30.864 28.628 47.792 28.716 ;
        RECT 47.332 12.16 110 15.5 ;
        RECT 47.746 11.746 47.792 28.716 ;
        RECT 30.818 28.674 47.746 28.762 ;
        RECT 47.378 12.114 110 15.5 ;
        RECT 47.7 11.792 47.746 28.762 ;
        RECT 30.772 28.72 47.7 28.808 ;
        RECT 47.424 12.068 110 15.5 ;
        RECT 47.654 11.838 47.7 28.808 ;
        RECT 30.726 28.766 47.654 28.854 ;
        RECT 47.47 12.022 110 15.5 ;
        RECT 47.608 11.884 47.654 28.854 ;
        RECT 30.68 28.812 47.608 28.9 ;
        RECT 47.516 11.976 110 15.5 ;
        RECT 47.562 11.93 47.608 28.9 ;
        RECT 30.634 28.858 47.562 28.946 ;
        RECT 30.588 28.904 47.516 28.992 ;
        RECT 30.542 28.95 47.47 29.038 ;
        RECT 30.496 28.996 47.424 29.084 ;
        RECT 30.45 29.042 47.378 29.13 ;
        RECT 30.404 29.088 47.332 29.176 ;
        RECT 30.358 29.134 47.286 29.222 ;
        RECT 30.312 29.18 47.24 29.268 ;
        RECT 30.266 29.226 47.194 29.314 ;
        RECT 30.22 29.272 47.148 29.36 ;
        RECT 30.174 29.318 47.102 29.406 ;
        RECT 30.128 29.364 47.056 29.452 ;
        RECT 30.082 29.41 47.01 29.498 ;
        RECT 30.036 29.456 46.964 29.544 ;
        RECT 29.99 29.502 46.918 29.59 ;
        RECT 29.944 29.548 46.872 29.636 ;
        RECT 29.898 29.594 46.826 29.682 ;
        RECT 29.852 29.64 46.78 29.728 ;
        RECT 29.806 29.686 46.734 29.774 ;
        RECT 29.76 29.732 46.688 29.82 ;
        RECT 29.714 29.778 46.642 29.866 ;
        RECT 29.668 29.824 46.596 29.912 ;
        RECT 29.622 29.87 46.55 29.958 ;
        RECT 29.576 29.916 46.504 30.004 ;
        RECT 29.53 29.962 46.458 30.05 ;
        RECT 29.484 30.008 46.412 30.096 ;
        RECT 29.438 30.054 46.366 30.142 ;
        RECT 29.392 30.1 46.32 30.188 ;
        RECT 29.346 30.146 46.274 30.234 ;
        RECT 29.3 30.192 46.228 30.28 ;
        RECT 29.254 30.238 46.182 30.326 ;
        RECT 29.208 30.284 46.136 30.372 ;
        RECT 29.162 30.33 46.09 30.418 ;
        RECT 29.116 30.376 46.044 30.464 ;
        RECT 29.07 30.422 45.998 30.51 ;
        RECT 29.024 30.468 45.952 30.556 ;
        RECT 28.978 30.514 45.906 30.602 ;
        RECT 28.932 30.56 45.86 30.648 ;
        RECT 28.886 30.606 45.814 30.694 ;
        RECT 28.84 30.652 45.768 30.74 ;
        RECT 28.794 30.698 45.722 30.786 ;
        RECT 28.748 30.744 45.676 30.832 ;
        RECT 28.702 30.79 45.63 30.878 ;
        RECT 28.656 30.836 45.584 30.924 ;
        RECT 28.61 30.882 45.538 30.97 ;
        RECT 28.564 30.928 45.492 31.016 ;
        RECT 28.518 30.974 45.446 31.062 ;
        RECT 28.472 31.02 45.4 31.108 ;
        RECT 28.426 31.066 45.354 31.154 ;
        RECT 28.38 31.112 45.308 31.2 ;
        RECT 28.334 31.158 45.262 31.246 ;
        RECT 28.288 31.204 45.216 31.292 ;
        RECT 28.242 31.25 45.17 31.338 ;
        RECT 28.196 31.296 45.124 31.384 ;
        RECT 28.15 31.342 45.078 31.43 ;
        RECT 28.104 31.388 45.032 31.476 ;
        RECT 28.058 31.434 44.986 31.522 ;
        RECT 28.012 31.48 44.94 31.568 ;
        RECT 27.966 31.526 44.894 31.614 ;
        RECT 27.92 31.572 44.848 31.66 ;
        RECT 27.874 31.618 44.802 31.706 ;
        RECT 27.828 31.664 44.756 31.752 ;
        RECT 27.782 31.71 44.71 31.798 ;
        RECT 27.736 31.756 44.664 31.844 ;
        RECT 27.69 31.802 44.618 31.89 ;
        RECT 27.644 31.848 44.572 31.936 ;
        RECT 27.598 31.894 44.526 31.982 ;
        RECT 27.552 31.94 44.48 32.028 ;
        RECT 27.506 31.986 44.434 32.074 ;
        RECT 27.46 32.032 44.388 32.12 ;
        RECT 27.414 32.078 44.342 32.166 ;
        RECT 27.368 32.124 44.296 32.212 ;
        RECT 27.322 32.17 44.25 32.258 ;
        RECT 27.276 32.216 44.204 32.304 ;
        RECT 27.23 32.262 44.158 32.35 ;
        RECT 27.184 32.308 44.112 32.396 ;
        RECT 27.138 32.354 44.066 32.442 ;
        RECT 27.092 32.4 44.02 32.488 ;
        RECT 27.046 32.446 43.974 32.534 ;
        RECT 27 32.492 43.928 32.58 ;
        RECT 26.954 32.538 43.882 32.626 ;
        RECT 26.908 32.584 43.836 32.672 ;
        RECT 26.862 32.63 43.79 32.718 ;
        RECT 26.816 32.676 43.744 32.764 ;
        RECT 26.77 32.722 43.698 32.81 ;
        RECT 26.724 32.768 43.652 32.856 ;
        RECT 26.678 32.814 43.606 32.902 ;
        RECT 26.632 32.86 43.56 32.948 ;
        RECT 26.586 32.906 43.514 32.994 ;
        RECT 26.54 32.952 43.468 33.04 ;
        RECT 26.494 32.998 43.422 33.086 ;
        RECT 26.448 33.044 43.376 33.132 ;
        RECT 26.402 33.09 43.33 33.178 ;
        RECT 26.356 33.136 43.284 33.224 ;
        RECT 26.31 33.182 43.238 33.27 ;
        RECT 26.264 33.228 43.192 33.316 ;
        RECT 26.218 33.274 43.146 33.362 ;
        RECT 26.172 33.32 43.1 33.408 ;
        RECT 26.126 33.366 43.054 33.454 ;
        RECT 26.08 33.412 43.008 33.5 ;
        RECT 26.034 33.458 42.962 33.546 ;
        RECT 25.988 33.504 42.916 33.592 ;
        RECT 25.942 33.55 42.87 33.638 ;
        RECT 25.896 33.596 42.824 33.684 ;
        RECT 25.85 33.642 42.778 33.73 ;
        RECT 25.804 33.688 42.732 33.776 ;
        RECT 25.758 33.734 42.686 33.822 ;
        RECT 25.712 33.78 42.64 33.868 ;
        RECT 25.666 33.826 42.594 33.914 ;
        RECT 25.62 33.872 42.548 33.96 ;
        RECT 25.574 33.918 42.502 34.006 ;
        RECT 25.528 33.964 42.456 34.052 ;
        RECT 25.482 34.01 42.41 34.098 ;
        RECT 25.436 34.056 42.364 34.144 ;
        RECT 25.39 34.102 42.318 34.19 ;
        RECT 25.344 34.148 42.272 34.236 ;
        RECT 25.298 34.194 42.226 34.282 ;
        RECT 25.252 34.24 42.18 34.328 ;
        RECT 25.206 34.286 42.134 34.374 ;
        RECT 25.16 34.332 42.088 34.42 ;
        RECT 25.114 34.378 42.042 34.466 ;
        RECT 25.068 34.424 41.996 34.512 ;
        RECT 25.022 34.47 41.95 34.558 ;
        RECT 24.976 34.516 41.904 34.604 ;
        RECT 24.93 34.562 41.858 34.65 ;
        RECT 24.884 34.608 41.812 34.696 ;
        RECT 24.838 34.654 41.766 34.742 ;
        RECT 24.792 34.7 41.72 34.788 ;
        RECT 24.746 34.746 41.674 34.834 ;
        RECT 24.7 34.792 41.628 34.88 ;
        RECT 24.654 34.838 41.582 34.926 ;
        RECT 24.608 34.884 41.536 34.972 ;
        RECT 24.562 34.93 41.49 35.018 ;
        RECT 24.516 34.976 41.444 35.064 ;
        RECT 24.47 35.022 41.398 35.11 ;
        RECT 24.424 35.068 41.352 35.156 ;
        RECT 24.378 35.114 41.306 35.202 ;
        RECT 24.332 35.16 41.26 35.248 ;
        RECT 24.286 35.206 41.214 35.294 ;
        RECT 24.24 35.252 41.168 35.34 ;
        RECT 24.194 35.298 41.122 35.386 ;
        RECT 24.148 35.344 41.076 35.432 ;
        RECT 24.102 35.39 41.03 35.478 ;
        RECT 24.056 35.436 40.984 35.524 ;
        RECT 24.01 35.482 40.938 35.57 ;
        RECT 23.964 35.528 40.892 35.616 ;
        RECT 23.918 35.574 40.846 35.662 ;
        RECT 23.872 35.62 40.8 35.708 ;
        RECT 23.826 35.666 40.754 35.754 ;
        RECT 23.78 35.712 40.708 35.8 ;
        RECT 23.734 35.758 40.662 35.846 ;
        RECT 23.688 35.804 40.616 35.892 ;
        RECT 23.642 35.85 40.57 35.938 ;
        RECT 23.596 35.896 40.524 35.984 ;
        RECT 23.55 35.942 40.478 36.03 ;
        RECT 23.504 35.988 40.432 36.076 ;
        RECT 23.458 36.034 40.386 36.122 ;
        RECT 23.412 36.08 40.34 36.168 ;
        RECT 23.366 36.126 40.294 36.214 ;
        RECT 23.32 36.172 40.248 36.26 ;
        RECT 23.274 36.218 40.202 36.306 ;
        RECT 23.228 36.264 40.156 36.352 ;
        RECT 23.182 36.31 40.11 36.398 ;
        RECT 23.136 36.356 40.064 36.444 ;
        RECT 23.09 36.402 40.018 36.49 ;
        RECT 23.044 36.448 39.972 36.536 ;
        RECT 22.998 36.494 39.926 36.582 ;
        RECT 22.952 36.54 39.88 36.628 ;
        RECT 22.906 36.586 39.834 36.674 ;
        RECT 22.86 36.632 39.788 36.72 ;
        RECT 22.814 36.678 39.742 36.766 ;
        RECT 22.768 36.724 39.696 36.812 ;
        RECT 22.722 36.77 39.65 36.858 ;
        RECT 22.676 36.816 39.604 36.904 ;
        RECT 22.63 36.862 39.558 36.95 ;
        RECT 22.584 36.908 39.512 36.996 ;
        RECT 22.538 36.954 39.466 37.042 ;
        RECT 22.492 37 39.42 37.088 ;
        RECT 22.446 37.046 39.374 37.134 ;
        RECT 22.4 37.092 39.328 37.18 ;
        RECT 22.354 37.138 39.282 37.226 ;
        RECT 22.308 37.184 39.236 37.272 ;
        RECT 22.262 37.23 39.19 37.318 ;
        RECT 22.216 37.276 39.144 37.364 ;
        RECT 22.17 37.322 39.098 37.41 ;
        RECT 22.124 37.368 39.052 37.456 ;
        RECT 22.078 37.414 39.006 37.502 ;
        RECT 22.032 37.46 38.96 37.548 ;
        RECT 21.986 37.506 38.914 37.594 ;
        RECT 21.94 37.552 38.868 37.64 ;
        RECT 21.894 37.598 38.822 37.686 ;
        RECT 21.848 37.644 38.776 37.732 ;
        RECT 21.802 37.69 38.73 37.778 ;
        RECT 21.756 37.736 38.684 37.824 ;
        RECT 21.71 37.782 38.638 37.87 ;
        RECT 21.664 37.828 38.592 37.916 ;
        RECT 21.618 37.874 38.546 37.962 ;
        RECT 21.572 37.92 38.5 38.008 ;
        RECT 21.526 37.966 38.454 38.054 ;
        RECT 21.48 38.012 38.408 38.1 ;
        RECT 21.434 38.058 38.362 38.146 ;
        RECT 21.388 38.104 38.316 38.192 ;
        RECT 21.342 38.15 38.27 38.238 ;
        RECT 21.296 38.196 38.224 38.284 ;
        RECT 21.25 38.242 38.178 38.33 ;
        RECT 21.204 38.288 38.132 38.376 ;
        RECT 21.158 38.334 38.086 38.422 ;
        RECT 21.112 38.38 38.04 38.468 ;
        RECT 21.066 38.426 37.994 38.514 ;
        RECT 21.02 38.472 37.948 38.56 ;
        RECT 20.974 38.518 37.902 38.606 ;
        RECT 20.928 38.564 37.856 38.652 ;
        RECT 20.882 38.61 37.81 38.698 ;
        RECT 20.836 38.656 37.764 38.744 ;
        RECT 20.79 38.702 37.718 38.79 ;
        RECT 20.744 38.748 37.672 38.836 ;
        RECT 20.698 38.794 37.626 38.882 ;
        RECT 20.652 38.84 37.58 38.928 ;
        RECT 20.606 38.886 37.534 38.974 ;
        RECT 20.56 38.932 37.488 39.02 ;
        RECT 20.514 38.978 37.442 39.066 ;
        RECT 20.468 39.024 37.396 39.112 ;
        RECT 20.422 39.07 37.35 39.158 ;
        RECT 20.376 39.116 37.304 39.204 ;
        RECT 20.33 39.162 37.258 39.25 ;
        RECT 20.284 39.208 37.212 39.296 ;
        RECT 20.238 39.254 37.166 39.342 ;
        RECT 20.192 39.3 37.12 39.388 ;
        RECT 20.146 39.346 37.074 39.434 ;
        RECT 20.1 39.392 37.028 39.48 ;
        RECT 20.054 39.438 36.982 39.526 ;
        RECT 20.008 39.484 36.936 39.572 ;
        RECT 19.962 39.53 36.89 39.618 ;
        RECT 19.916 39.576 36.844 39.664 ;
        RECT 19.87 39.622 36.798 39.71 ;
        RECT 19.824 39.668 36.752 39.756 ;
        RECT 19.778 39.714 36.706 39.802 ;
        RECT 19.732 39.76 36.66 39.848 ;
        RECT 19.686 39.806 36.614 39.894 ;
        RECT 19.64 39.852 36.568 39.94 ;
        RECT 19.594 39.898 36.522 39.986 ;
        RECT 19.548 39.944 36.476 40.032 ;
        RECT 19.502 39.99 36.43 40.078 ;
        RECT 19.456 40.036 36.384 40.124 ;
        RECT 19.41 40.082 36.338 40.17 ;
        RECT 19.364 40.128 36.292 40.216 ;
        RECT 19.318 40.174 36.246 40.262 ;
        RECT 19.272 40.22 36.2 40.308 ;
        RECT 19.226 40.266 36.154 40.354 ;
        RECT 19.18 40.312 36.108 40.4 ;
        RECT 19.134 40.358 36.062 40.446 ;
        RECT 19.088 40.404 36.016 40.492 ;
        RECT 19.042 40.45 35.97 40.538 ;
        RECT 18.996 40.496 35.924 40.584 ;
        RECT 18.95 40.542 35.878 40.63 ;
        RECT 18.904 40.588 35.832 40.676 ;
        RECT 18.858 40.634 35.786 40.722 ;
        RECT 18.812 40.68 35.74 40.768 ;
        RECT 18.766 40.726 35.694 40.814 ;
        RECT 18.72 40.772 35.648 40.86 ;
        RECT 18.674 40.818 35.602 40.906 ;
        RECT 18.628 40.864 35.556 40.952 ;
        RECT 18.582 40.91 35.51 40.998 ;
        RECT 18.536 40.956 35.464 41.044 ;
        RECT 18.49 41.002 35.418 41.09 ;
        RECT 18.444 41.048 35.372 41.136 ;
        RECT 18.398 41.094 35.326 41.182 ;
        RECT 18.352 41.14 35.28 41.228 ;
        RECT 18.306 41.186 35.234 41.274 ;
        RECT 18.26 41.232 35.188 41.32 ;
        RECT 18.214 41.278 35.142 41.366 ;
        RECT 18.168 41.324 35.096 41.412 ;
        RECT 18.122 41.37 35.05 41.458 ;
        RECT 18.076 41.416 35.004 41.504 ;
        RECT 18.03 41.462 34.958 41.55 ;
        RECT 17.984 41.508 34.912 41.596 ;
        RECT 17.938 41.554 34.866 41.642 ;
        RECT 17.892 41.6 34.82 41.688 ;
        RECT 17.846 41.646 34.774 41.734 ;
        RECT 17.8 41.692 34.728 41.78 ;
        RECT 17.754 41.738 34.682 41.826 ;
        RECT 17.708 41.784 34.636 41.872 ;
        RECT 17.662 41.83 34.59 41.918 ;
        RECT 17.616 41.876 34.544 41.964 ;
        RECT 17.57 41.922 34.498 42.01 ;
        RECT 17.524 41.968 34.452 42.056 ;
        RECT 17.478 42.014 34.406 42.102 ;
        RECT 17.432 42.06 34.36 42.148 ;
        RECT 17.386 42.106 34.314 42.194 ;
        RECT 17.34 42.152 34.268 42.24 ;
        RECT 17.294 42.198 34.222 42.286 ;
        RECT 17.248 42.244 34.176 42.332 ;
        RECT 17.202 42.29 34.13 42.378 ;
        RECT 17.156 42.336 34.084 42.424 ;
        RECT 17.11 42.382 34.038 42.47 ;
        RECT 17.064 42.428 33.992 42.516 ;
        RECT 17.018 42.474 33.946 42.562 ;
        RECT 16.972 42.52 33.9 42.608 ;
        RECT 16.926 42.566 33.854 42.654 ;
        RECT 16.88 42.612 33.808 42.7 ;
        RECT 16.834 42.658 33.762 42.746 ;
        RECT 16.788 42.704 33.716 42.792 ;
        RECT 16.742 42.75 33.67 42.838 ;
        RECT 16.696 42.796 33.624 42.884 ;
        RECT 16.65 42.842 33.578 42.93 ;
        RECT 16.604 42.888 33.532 42.976 ;
        RECT 16.558 42.934 33.486 43.022 ;
        RECT 16.512 42.98 33.44 43.068 ;
        RECT 16.466 43.026 33.394 43.114 ;
        RECT 16.42 43.072 33.348 43.16 ;
        RECT 16.374 43.118 33.302 43.206 ;
        RECT 16.328 43.164 33.256 43.252 ;
        RECT 16.282 43.21 33.21 43.298 ;
        RECT 16.236 43.256 33.164 43.344 ;
        RECT 16.19 43.302 33.118 43.39 ;
        RECT 16.144 43.348 33.072 43.436 ;
        RECT 16.098 43.394 33.026 43.482 ;
        RECT 16.052 43.44 32.98 43.528 ;
        RECT 16.006 43.486 32.934 43.574 ;
        RECT 15.96 43.532 32.888 43.62 ;
        RECT 15.914 43.578 32.842 43.666 ;
        RECT 15.868 43.624 32.796 43.712 ;
        RECT 15.822 43.67 32.75 43.758 ;
        RECT 15.776 43.716 32.704 43.804 ;
        RECT 15.73 43.762 32.658 43.85 ;
        RECT 15.684 43.808 32.612 43.896 ;
        RECT 15.638 43.854 32.566 43.942 ;
        RECT 15.592 43.9 32.52 43.988 ;
        RECT 15.5 43.992 32.474 44.034 ;
        RECT 15.546 43.946 32.474 44.034 ;
        RECT 15.46 44.035 32.428 44.08 ;
        RECT 15.414 44.078 32.382 44.126 ;
        RECT 15.368 44.124 32.336 44.172 ;
        RECT 15.322 44.17 32.29 44.218 ;
        RECT 15.276 44.216 32.244 44.264 ;
        RECT 15.23 44.262 32.198 44.31 ;
        RECT 15.184 44.308 32.152 44.356 ;
        RECT 15.138 44.354 32.106 44.402 ;
        RECT 15.092 44.4 32.06 44.448 ;
        RECT 15.046 44.446 32.014 44.494 ;
        RECT 15 44.492 31.968 44.54 ;
        RECT 14.954 44.538 31.922 44.586 ;
        RECT 14.908 44.584 31.876 44.632 ;
        RECT 14.862 44.63 31.83 44.678 ;
        RECT 14.816 44.676 31.784 44.724 ;
        RECT 14.77 44.722 31.738 44.77 ;
        RECT 14.724 44.768 31.692 44.816 ;
        RECT 14.678 44.814 31.646 44.862 ;
        RECT 14.632 44.86 31.6 44.908 ;
        RECT 14.586 44.906 31.554 44.954 ;
        RECT 14.54 44.952 31.508 45 ;
        RECT 14.494 44.998 31.462 45.046 ;
        RECT 14.448 45.044 31.416 45.092 ;
        RECT 14.402 45.09 31.37 45.138 ;
        RECT 14.356 45.136 31.324 45.184 ;
        RECT 14.31 45.182 31.278 45.23 ;
        RECT 14.264 45.228 31.232 45.276 ;
        RECT 14.218 45.274 31.186 45.322 ;
        RECT 14.172 45.32 31.14 45.368 ;
        RECT 14.126 45.366 31.094 45.414 ;
        RECT 14.08 45.412 31.048 45.46 ;
        RECT 14.034 45.458 31.002 45.506 ;
        RECT 13.988 45.504 30.956 45.552 ;
        RECT 13.942 45.55 30.91 45.598 ;
        RECT 13.896 45.596 30.864 45.644 ;
        RECT 13.85 45.642 30.818 45.69 ;
        RECT 13.804 45.688 30.772 45.736 ;
        RECT 13.758 45.734 30.726 45.782 ;
        RECT 13.712 45.78 30.68 45.828 ;
        RECT 13.666 45.826 30.634 45.874 ;
        RECT 13.62 45.872 30.588 45.92 ;
        RECT 13.574 45.918 30.542 45.966 ;
        RECT 13.528 45.964 30.496 46.012 ;
        RECT 13.482 46.01 30.45 46.058 ;
        RECT 13.436 46.056 30.404 46.104 ;
        RECT 13.39 46.102 30.358 46.15 ;
        RECT 13.344 46.148 30.312 46.196 ;
        RECT 13.298 46.194 30.266 46.242 ;
        RECT 13.252 46.24 30.22 46.288 ;
        RECT 13.206 46.286 30.174 46.334 ;
        RECT 13.16 46.332 30.128 46.38 ;
        RECT 13.114 46.378 30.082 46.426 ;
        RECT 13.068 46.424 30.036 46.472 ;
        RECT 13.022 46.47 29.99 46.518 ;
        RECT 12.976 46.516 29.944 46.564 ;
        RECT 12.93 46.562 29.898 46.61 ;
        RECT 12.884 46.608 29.852 46.656 ;
        RECT 12.838 46.654 29.806 46.702 ;
        RECT 12.792 46.7 29.76 46.748 ;
        RECT 12.746 46.746 29.714 46.794 ;
        RECT 12.7 46.792 29.668 46.84 ;
        RECT 12.654 46.838 29.622 46.886 ;
        RECT 12.608 46.884 29.576 46.932 ;
        RECT 12.562 46.93 29.53 46.978 ;
        RECT 12.516 46.976 29.484 47.024 ;
        RECT 12.47 47.022 29.438 47.07 ;
        RECT 12.424 47.068 29.392 47.116 ;
        RECT 12.378 47.114 29.346 47.162 ;
        RECT 12.332 47.16 29.3 47.208 ;
        RECT 12.286 47.206 29.254 47.254 ;
        RECT 12.24 47.252 29.208 47.3 ;
        RECT 12.194 47.298 29.162 47.346 ;
        RECT 12.148 47.344 29.116 47.392 ;
        RECT 12.102 47.39 29.07 47.438 ;
        RECT 12.056 47.436 29.024 47.484 ;
        RECT 12.01 47.482 28.978 47.53 ;
        RECT 11.964 47.528 28.932 47.576 ;
        RECT 11.918 47.574 28.886 47.622 ;
        RECT 11.872 47.62 28.84 47.668 ;
        RECT 11.826 47.666 28.794 47.714 ;
        RECT 11.78 47.712 28.748 47.76 ;
        RECT 11.734 47.758 28.702 47.806 ;
        RECT 11.688 47.804 28.656 47.852 ;
        RECT 11.642 47.85 28.61 47.898 ;
        RECT 11.596 47.896 28.564 47.944 ;
        RECT 11.55 47.942 28.518 47.99 ;
        RECT 11.504 47.988 28.472 48.036 ;
        RECT 11.458 48.034 28.426 48.082 ;
        RECT 11.412 48.08 28.38 48.128 ;
        RECT 11.366 48.126 28.334 48.174 ;
        RECT 11.32 48.172 28.288 48.22 ;
        RECT 11.274 48.218 28.242 48.266 ;
        RECT 11.228 48.264 28.196 48.312 ;
        RECT 11.182 48.31 28.15 48.358 ;
        RECT 11.136 48.356 28.104 48.404 ;
        RECT 11.09 48.402 28.058 48.45 ;
        RECT 11.044 48.448 28.012 48.496 ;
        RECT 10.998 48.494 27.966 48.542 ;
        RECT 10.952 48.54 27.92 48.588 ;
        RECT 10.906 48.586 27.874 48.634 ;
        RECT 10.86 48.632 27.828 48.68 ;
        RECT 10.814 48.678 27.782 48.726 ;
        RECT 10.768 48.724 27.736 48.772 ;
        RECT 10.722 48.77 27.69 48.818 ;
        RECT 10.676 48.816 27.644 48.864 ;
        RECT 10.63 48.862 27.598 48.91 ;
        RECT 10.584 48.908 27.552 48.956 ;
        RECT 10.538 48.954 27.506 49.002 ;
        RECT 10.492 49 27.46 49.048 ;
        RECT 10.446 49.046 27.414 49.094 ;
        RECT 10.4 49.092 27.368 49.14 ;
        RECT 10.354 49.138 27.322 49.186 ;
        RECT 10.308 49.184 27.276 49.232 ;
        RECT 10.262 49.23 27.23 49.278 ;
        RECT 10.216 49.276 27.184 49.324 ;
        RECT 10.17 49.322 27.138 49.37 ;
        RECT 10.124 49.368 27.092 49.416 ;
        RECT 10.078 49.414 27.046 49.462 ;
      LAYER MET2 ;
        RECT 28.362 51.38 45.33 51.428 ;
        RECT 28.316 51.426 45.284 51.474 ;
        RECT 28.27 51.472 45.238 51.52 ;
        RECT 28.224 51.518 45.192 51.566 ;
        RECT 28.178 51.564 45.146 51.612 ;
        RECT 28.132 51.61 45.1 51.658 ;
        RECT 28.086 51.656 45.054 51.704 ;
        RECT 28.04 51.702 45.008 51.75 ;
        RECT 27.994 51.748 44.962 51.796 ;
        RECT 27.948 51.794 44.916 51.842 ;
        RECT 27.902 51.84 44.87 51.888 ;
        RECT 27.856 51.886 44.824 51.934 ;
        RECT 27.81 51.932 44.778 51.98 ;
        RECT 27.764 51.978 44.732 52.026 ;
        RECT 27.718 52.024 44.686 52.072 ;
        RECT 27.672 52.07 44.64 52.118 ;
        RECT 27.626 52.116 44.594 52.164 ;
        RECT 27.58 52.162 44.548 52.21 ;
        RECT 27.534 52.208 44.502 52.256 ;
        RECT 27.488 52.254 44.456 52.302 ;
        RECT 27.442 52.3 44.41 52.348 ;
        RECT 27.396 52.346 44.364 52.394 ;
        RECT 27.35 52.392 44.318 52.44 ;
        RECT 27.304 52.438 44.272 52.486 ;
        RECT 27.258 52.484 44.226 52.532 ;
        RECT 27.212 52.53 44.18 52.578 ;
        RECT 27.166 52.576 44.134 52.624 ;
        RECT 27.12 52.622 44.088 52.67 ;
        RECT 27.074 52.668 44.042 52.716 ;
        RECT 27.028 52.714 43.996 52.762 ;
        RECT 26.982 52.76 43.95 52.808 ;
        RECT 26.936 52.806 43.904 52.854 ;
        RECT 26.89 52.852 43.858 52.9 ;
        RECT 26.844 52.898 43.812 52.946 ;
        RECT 26.798 52.944 43.766 52.992 ;
        RECT 26.752 52.99 43.72 53.038 ;
        RECT 26.706 53.036 43.674 53.084 ;
        RECT 26.66 53.082 43.628 53.13 ;
        RECT 26.614 53.128 43.582 53.176 ;
        RECT 26.568 53.174 43.536 53.222 ;
        RECT 26.522 53.22 43.49 53.268 ;
        RECT 26.476 53.266 43.444 53.314 ;
        RECT 26.43 53.312 43.398 53.36 ;
        RECT 26.384 53.358 43.352 53.406 ;
        RECT 26.338 53.404 43.306 53.452 ;
        RECT 26.292 53.45 43.26 53.498 ;
        RECT 26.246 53.496 43.214 53.544 ;
        RECT 26.2 53.542 43.168 53.59 ;
        RECT 26.154 53.588 43.122 53.636 ;
        RECT 26.108 53.634 43.076 53.682 ;
        RECT 26.062 53.68 43.03 53.728 ;
        RECT 26.016 53.726 42.984 53.774 ;
        RECT 25.97 53.772 42.938 53.82 ;
        RECT 25.924 53.818 42.892 53.866 ;
        RECT 25.878 53.864 42.846 53.912 ;
        RECT 25.832 53.91 42.8 53.958 ;
        RECT 25.786 53.956 42.754 54.004 ;
        RECT 25.74 54.002 42.708 54.05 ;
        RECT 25.694 54.048 42.662 54.096 ;
        RECT 25.648 54.094 42.616 54.142 ;
        RECT 25.602 54.14 42.57 54.188 ;
        RECT 25.556 54.186 42.524 54.234 ;
        RECT 25.51 54.232 42.478 54.28 ;
        RECT 25.464 54.278 42.432 54.326 ;
        RECT 25.418 54.324 42.386 54.372 ;
        RECT 25.372 54.37 42.34 54.418 ;
        RECT 25.326 54.416 42.294 54.464 ;
        RECT 25.28 54.462 42.248 54.51 ;
        RECT 25.234 54.508 42.202 54.556 ;
        RECT 25.188 54.554 42.156 54.602 ;
        RECT 25.142 54.6 42.11 54.648 ;
        RECT 25.096 54.646 42.064 54.694 ;
        RECT 25.05 54.692 42.018 54.74 ;
        RECT 25.004 54.738 41.972 54.786 ;
        RECT 24.958 54.784 41.926 54.832 ;
        RECT 24.912 54.83 41.88 54.878 ;
        RECT 24.866 54.876 41.834 54.924 ;
        RECT 24.82 54.922 41.788 54.97 ;
        RECT 24.774 54.968 41.742 55.016 ;
        RECT 24.728 55.014 41.696 55.062 ;
        RECT 24.682 55.06 41.65 55.108 ;
        RECT 24.636 55.106 41.604 55.154 ;
        RECT 24.59 55.152 41.558 55.2 ;
        RECT 24.544 55.198 41.512 55.246 ;
        RECT 24.498 55.244 41.466 55.292 ;
        RECT 24.452 55.29 41.42 55.338 ;
        RECT 24.406 55.336 41.374 55.384 ;
        RECT 24.36 55.382 41.328 55.43 ;
        RECT 24.314 55.428 41.282 55.476 ;
        RECT 24.268 55.474 41.236 55.522 ;
        RECT 24.222 55.52 41.19 55.568 ;
        RECT 24.176 55.566 41.144 55.614 ;
        RECT 24.13 55.612 41.098 55.66 ;
        RECT 24.084 55.658 41.052 55.706 ;
        RECT 24.038 55.704 41.006 55.752 ;
        RECT 23.992 55.75 40.96 55.798 ;
        RECT 23.946 55.796 40.914 55.844 ;
        RECT 23.9 55.842 40.868 55.89 ;
        RECT 23.854 55.888 40.822 55.936 ;
        RECT 23.808 55.934 40.776 55.982 ;
        RECT 23.762 55.98 40.73 56.028 ;
        RECT 23.716 56.026 40.684 56.074 ;
        RECT 23.67 56.072 40.638 56.12 ;
        RECT 23.624 56.118 40.592 56.166 ;
        RECT 23.578 56.164 40.546 56.212 ;
        RECT 23.532 56.21 40.5 56.258 ;
        RECT 23.486 56.256 40.454 56.304 ;
        RECT 23.44 56.302 40.408 56.35 ;
        RECT 23.394 56.348 40.362 56.396 ;
        RECT 23.348 56.394 40.316 56.442 ;
        RECT 23.302 56.44 40.27 56.488 ;
        RECT 23.256 56.486 40.224 56.534 ;
        RECT 23.21 56.532 40.178 56.58 ;
        RECT 23.164 56.578 40.132 56.626 ;
        RECT 23.118 56.624 40.086 56.672 ;
        RECT 23.072 56.67 40.04 56.718 ;
        RECT 23.026 56.716 39.994 56.764 ;
        RECT 22.98 56.762 39.948 56.81 ;
        RECT 22.934 56.808 39.902 56.856 ;
        RECT 22.888 56.854 39.856 56.902 ;
        RECT 22.842 56.9 39.81 56.948 ;
        RECT 22.796 56.946 39.764 56.994 ;
        RECT 22.75 56.992 39.718 57.04 ;
        RECT 22.704 57.038 39.672 57.086 ;
        RECT 22.658 57.084 39.626 57.132 ;
        RECT 22.612 57.13 39.58 57.178 ;
        RECT 22.566 57.176 39.534 57.224 ;
        RECT 22.52 57.222 39.488 57.27 ;
        RECT 22.474 57.268 39.442 57.316 ;
        RECT 22.428 57.314 39.396 57.362 ;
        RECT 22.382 57.36 39.35 57.408 ;
        RECT 22.336 57.406 39.304 57.454 ;
        RECT 22.29 57.452 39.258 57.5 ;
        RECT 22.244 57.498 39.212 57.546 ;
        RECT 22.198 57.544 39.166 57.592 ;
        RECT 22.152 57.59 39.12 57.638 ;
        RECT 22.106 57.636 39.074 57.684 ;
        RECT 22.06 57.682 39.028 57.73 ;
        RECT 22.014 57.728 38.982 57.776 ;
        RECT 21.968 57.774 38.936 57.822 ;
        RECT 21.922 57.82 38.89 57.868 ;
        RECT 21.876 57.866 38.844 57.914 ;
        RECT 21.83 57.912 38.798 57.96 ;
        RECT 21.784 57.958 38.752 58.006 ;
        RECT 21.738 58.004 38.706 58.052 ;
        RECT 21.692 58.05 38.66 58.098 ;
        RECT 21.646 58.096 38.614 58.144 ;
        RECT 21.6 58.142 38.568 58.19 ;
        RECT 21.554 58.188 38.522 58.236 ;
        RECT 21.508 58.234 38.476 58.282 ;
        RECT 21.462 58.28 38.43 58.328 ;
        RECT 21.416 58.326 38.384 58.374 ;
        RECT 21.37 58.372 38.338 58.42 ;
        RECT 21.324 58.418 38.292 58.466 ;
        RECT 21.278 58.464 38.246 58.512 ;
        RECT 21.232 58.51 38.2 58.558 ;
        RECT 21.186 58.556 38.154 58.604 ;
        RECT 21.14 58.602 38.108 58.65 ;
        RECT 21.094 58.648 38.062 58.696 ;
        RECT 21.048 58.694 38.016 58.742 ;
        RECT 21.002 58.74 37.97 58.788 ;
        RECT 20.956 58.786 37.924 58.834 ;
        RECT 20.91 58.832 37.878 58.88 ;
        RECT 20.864 58.878 37.832 58.926 ;
        RECT 20.818 58.924 37.786 58.972 ;
        RECT 20.772 58.97 37.74 59.018 ;
        RECT 20.726 59.016 37.694 59.064 ;
        RECT 20.68 59.062 37.648 59.11 ;
        RECT 20.634 59.108 37.602 59.156 ;
        RECT 20.588 59.154 37.556 59.202 ;
        RECT 20.542 59.2 37.51 59.248 ;
        RECT 20.496 59.246 37.464 59.294 ;
        RECT 20.45 59.292 37.418 59.34 ;
        RECT 20.404 59.338 37.372 59.386 ;
        RECT 20.358 59.384 37.326 59.432 ;
        RECT 20.312 59.43 37.28 59.478 ;
        RECT 20.266 59.476 37.234 59.524 ;
        RECT 20.22 59.522 37.188 59.57 ;
        RECT 20.174 59.568 37.142 59.616 ;
        RECT 20.128 59.614 37.096 59.662 ;
        RECT 20.082 59.66 37.05 59.708 ;
        RECT 20.036 59.706 37.004 59.754 ;
        RECT 19.99 59.752 36.958 59.8 ;
        RECT 19.944 59.798 36.912 59.846 ;
        RECT 19.898 59.844 36.866 59.892 ;
        RECT 19.852 59.89 36.82 59.938 ;
        RECT 19.806 59.936 36.774 59.984 ;
        RECT 19.76 59.982 36.728 60.03 ;
        RECT 19.714 60.028 36.682 60.076 ;
        RECT 19.668 60.074 36.636 60.122 ;
        RECT 19.622 60.12 36.59 60.168 ;
        RECT 19.576 60.166 36.544 60.214 ;
        RECT 19.53 60.212 36.498 60.26 ;
        RECT 19.484 60.258 36.452 60.306 ;
        RECT 19.438 60.304 36.406 60.352 ;
        RECT 19.392 60.35 36.36 60.398 ;
        RECT 19.346 60.396 36.314 60.444 ;
        RECT 19.3 60.442 36.268 60.49 ;
        RECT 19.254 60.488 36.222 60.536 ;
        RECT 19.208 60.534 36.176 60.582 ;
        RECT 19.162 60.58 36.13 60.628 ;
        RECT 19.116 60.626 36.084 60.674 ;
        RECT 19.07 60.672 36.038 60.72 ;
        RECT 19.024 60.718 35.992 60.766 ;
        RECT 18.978 60.764 35.946 60.812 ;
        RECT 18.932 60.81 35.9 60.858 ;
        RECT 18.886 60.856 35.854 60.904 ;
        RECT 18.84 60.902 35.808 60.95 ;
        RECT 18.794 60.948 35.762 60.996 ;
        RECT 18.748 60.994 35.716 61.042 ;
        RECT 18.702 61.04 35.67 61.088 ;
        RECT 18.656 61.086 35.624 61.134 ;
        RECT 18.61 61.132 35.578 61.18 ;
        RECT 18.564 61.178 35.532 61.226 ;
        RECT 18.518 61.224 35.486 61.272 ;
        RECT 18.472 61.27 35.44 61.318 ;
        RECT 18.426 61.316 35.394 61.364 ;
        RECT 18.38 61.362 35.348 61.41 ;
        RECT 18.334 61.408 35.302 61.456 ;
        RECT 18.288 61.454 35.256 61.502 ;
        RECT 18.242 61.5 35.21 61.548 ;
        RECT 18.196 61.546 35.164 61.594 ;
        RECT 18.15 61.592 35.118 61.64 ;
        RECT 18.104 61.638 35.072 61.686 ;
        RECT 18.058 61.684 35.026 61.732 ;
        RECT 18.012 61.73 34.98 61.778 ;
        RECT 17.966 61.776 34.934 61.824 ;
        RECT 17.92 61.822 34.888 61.87 ;
        RECT 17.874 61.868 34.842 61.916 ;
        RECT 17.828 61.914 34.796 61.962 ;
        RECT 17.782 61.96 34.75 62.008 ;
        RECT 17.736 62.006 34.704 62.054 ;
        RECT 17.69 62.052 34.658 62.1 ;
        RECT 17.644 62.098 34.612 62.146 ;
        RECT 17.598 62.144 34.566 62.192 ;
        RECT 17.552 62.19 34.52 62.238 ;
        RECT 17.506 62.236 34.474 62.284 ;
        RECT 17.46 62.282 34.428 62.33 ;
        RECT 17.414 62.328 34.382 62.376 ;
        RECT 17.368 62.374 34.336 62.422 ;
        RECT 17.322 62.42 34.29 62.468 ;
        RECT 17.276 62.466 34.244 62.514 ;
        RECT 17.23 62.512 34.198 62.56 ;
        RECT 17.184 62.558 34.152 62.606 ;
        RECT 17.138 62.604 34.106 62.652 ;
        RECT 17.092 62.65 34.06 62.698 ;
        RECT 17.046 62.696 34.014 62.744 ;
        RECT 17 62.742 33.968 62.79 ;
        RECT 17 62.742 33.922 62.836 ;
        RECT 17 62.742 33.876 62.882 ;
        RECT 17 62.742 33.83 62.928 ;
        RECT 17 62.742 33.784 62.974 ;
        RECT 17 62.742 33.738 63.02 ;
        RECT 17 62.742 33.692 63.066 ;
        RECT 17 62.742 33.646 63.112 ;
        RECT 17 62.742 33.6 63.158 ;
        RECT 17 62.742 33.554 63.204 ;
        RECT 17 62.742 33.508 63.25 ;
        RECT 17 62.742 33.462 63.296 ;
        RECT 17 62.742 33.416 63.342 ;
        RECT 17 62.742 33.37 63.388 ;
        RECT 17 62.742 33.324 63.434 ;
        RECT 17 62.742 33.278 63.48 ;
        RECT 17 62.742 33.232 63.526 ;
        RECT 17 62.742 33.186 63.572 ;
        RECT 17 62.742 33.14 63.618 ;
        RECT 17 62.742 33.094 63.664 ;
        RECT 17 62.742 33.048 63.71 ;
        RECT 17 62.742 33.002 63.756 ;
        RECT 17 62.742 32.956 63.802 ;
        RECT 17 62.742 32.91 63.848 ;
        RECT 17 62.742 32.864 63.894 ;
        RECT 17 62.742 32.818 63.94 ;
        RECT 17 62.742 32.772 63.986 ;
        RECT 17 62.742 32.726 64.032 ;
        RECT 17 62.742 32.68 64.078 ;
        RECT 17 62.742 32.634 64.124 ;
        RECT 17 62.742 32.588 64.17 ;
        RECT 17 62.742 32.542 64.216 ;
        RECT 17 62.742 32.496 64.262 ;
        RECT 17 62.742 32.45 64.308 ;
        RECT 17 62.742 32.404 64.354 ;
        RECT 17 62.742 32.358 64.4 ;
        RECT 17 62.742 32.312 64.446 ;
        RECT 17 62.742 32.266 64.492 ;
        RECT 17 62.742 32.22 64.538 ;
        RECT 17 62.742 32.174 64.584 ;
        RECT 17 62.742 32.128 64.63 ;
        RECT 17 62.742 32.082 64.676 ;
        RECT 17 62.742 32.036 64.722 ;
        RECT 17 62.742 31.99 64.768 ;
        RECT 17 62.742 31.944 64.814 ;
        RECT 17 62.742 31.898 64.86 ;
        RECT 17 62.742 31.852 64.906 ;
        RECT 17 62.742 31.806 64.952 ;
        RECT 17 62.742 31.76 64.998 ;
        RECT 17 62.742 31.714 65.044 ;
        RECT 17 62.742 31.668 65.09 ;
        RECT 17 62.742 31.622 65.136 ;
        RECT 17 62.742 31.576 65.182 ;
        RECT 17 62.742 31.53 65.228 ;
        RECT 17 62.742 31.484 65.274 ;
        RECT 17 62.742 31.438 65.32 ;
        RECT 17 62.742 31.392 65.366 ;
        RECT 17 62.742 31.346 65.412 ;
        RECT 17 62.742 31.3 65.458 ;
        RECT 17 62.742 31.254 65.504 ;
        RECT 17 62.742 31.208 65.55 ;
        RECT 17 62.742 31.162 65.596 ;
        RECT 17 62.742 31.116 65.642 ;
        RECT 17 62.742 31.07 65.688 ;
        RECT 17 62.742 31.024 65.734 ;
        RECT 17 62.742 30.978 65.78 ;
        RECT 17 62.742 30.932 65.826 ;
        RECT 17 62.742 30.886 65.872 ;
        RECT 17 62.742 30.84 65.918 ;
        RECT 17 62.742 30.794 65.964 ;
        RECT 17 62.742 30.748 66.01 ;
        RECT 17 62.742 30.702 66.056 ;
        RECT 17 62.742 30.656 66.102 ;
        RECT 17 62.742 30.61 66.148 ;
        RECT 17 62.742 30.564 66.194 ;
        RECT 17 62.742 30.518 66.24 ;
        RECT 17 62.742 30.472 66.286 ;
        RECT 17 62.742 30.426 66.332 ;
        RECT 17 62.742 30.38 66.378 ;
        RECT 17 62.742 30.334 66.424 ;
        RECT 17 62.742 30.288 66.47 ;
        RECT 17 62.742 30.242 66.516 ;
        RECT 17 62.742 30.196 66.562 ;
        RECT 17 62.742 30.15 66.608 ;
        RECT 17 62.742 30.104 66.654 ;
        RECT 17 62.742 30.058 66.7 ;
        RECT 17 62.742 30.012 66.746 ;
        RECT 17 62.742 29.966 66.792 ;
        RECT 17 62.742 29.92 66.838 ;
        RECT 17 62.742 29.874 66.884 ;
        RECT 17 62.742 29.828 66.93 ;
        RECT 17 62.742 29.782 66.976 ;
        RECT 17 62.742 29.736 67.022 ;
        RECT 17 62.742 29.69 67.068 ;
        RECT 17 62.742 29.644 67.114 ;
        RECT 17 62.742 29.598 67.16 ;
        RECT 17 62.742 29.552 67.206 ;
        RECT 17 62.742 29.506 67.252 ;
        RECT 17 62.742 29.46 67.298 ;
        RECT 17 62.742 29.414 67.344 ;
        RECT 17 62.742 29.368 67.39 ;
        RECT 17 62.742 29.322 67.436 ;
        RECT 17 62.742 29.276 67.482 ;
        RECT 17 62.742 29.23 67.528 ;
        RECT 17 62.742 29.184 67.574 ;
        RECT 17 62.742 29.138 67.62 ;
        RECT 17 62.742 29.092 67.666 ;
        RECT 17 62.742 29.046 67.712 ;
        RECT 17 62.742 29 110 ;
        RECT 92.47 78.5 110 89.5 ;
        RECT 81.444 89.503 97.024 89.529 ;
        RECT 78.5 92.447 94.034 92.519 ;
        RECT 78.5 92.447 93.988 92.565 ;
        RECT 78.5 92.447 93.942 92.611 ;
        RECT 78.5 92.447 93.896 92.657 ;
        RECT 78.5 92.447 93.85 92.703 ;
        RECT 78.5 92.447 93.804 92.749 ;
        RECT 78.5 92.447 93.758 92.795 ;
        RECT 78.5 92.447 93.712 92.841 ;
        RECT 78.5 92.447 93.666 92.887 ;
        RECT 78.5 92.447 93.62 92.933 ;
        RECT 78.5 92.447 93.574 92.979 ;
        RECT 78.5 92.447 93.528 93.025 ;
        RECT 78.5 92.447 93.482 93.071 ;
        RECT 78.5 92.447 93.436 93.117 ;
        RECT 78.5 92.447 93.39 93.163 ;
        RECT 78.5 92.447 93.344 93.209 ;
        RECT 78.5 92.447 93.298 93.255 ;
        RECT 78.5 92.447 93.252 93.301 ;
        RECT 78.5 92.447 93.206 93.347 ;
        RECT 78.5 92.447 93.16 93.393 ;
        RECT 78.5 92.447 93.114 93.439 ;
        RECT 78.5 92.447 93.068 93.485 ;
        RECT 78.5 92.447 93.022 93.531 ;
        RECT 78.5 92.447 92.976 93.577 ;
        RECT 78.5 92.447 92.93 93.623 ;
        RECT 78.5 92.447 92.884 93.669 ;
        RECT 78.5 92.447 92.838 93.715 ;
        RECT 78.5 92.447 92.792 93.761 ;
        RECT 78.5 92.447 92.746 93.807 ;
        RECT 78.5 92.447 92.7 93.853 ;
        RECT 78.5 92.447 92.654 93.899 ;
        RECT 78.5 92.447 92.608 93.945 ;
        RECT 78.5 92.447 92.562 93.991 ;
        RECT 78.5 92.447 92.516 94.037 ;
        RECT 78.546 92.401 94.08 92.473 ;
        RECT 92.444 78.513 92.47 94.073 ;
        RECT 78.592 92.355 94.126 92.427 ;
        RECT 92.398 78.549 92.444 94.109 ;
        RECT 78.638 92.309 94.172 92.381 ;
        RECT 92.352 78.595 92.398 94.155 ;
        RECT 78.684 92.263 94.218 92.335 ;
        RECT 92.306 78.641 92.352 94.201 ;
        RECT 78.73 92.217 94.264 92.289 ;
        RECT 92.26 78.687 92.306 94.247 ;
        RECT 78.776 92.171 94.31 92.243 ;
        RECT 92.214 78.733 92.26 94.293 ;
        RECT 78.822 92.125 94.356 92.197 ;
        RECT 92.168 78.779 92.214 94.339 ;
        RECT 78.868 92.079 94.402 92.151 ;
        RECT 92.122 78.825 92.168 94.385 ;
        RECT 78.914 92.033 94.448 92.105 ;
        RECT 92.076 78.871 92.122 94.431 ;
        RECT 78.96 91.987 94.494 92.059 ;
        RECT 92.03 78.917 92.076 94.477 ;
        RECT 79.006 91.941 94.54 92.013 ;
        RECT 91.984 78.963 92.03 94.523 ;
        RECT 79.052 91.895 94.586 91.967 ;
        RECT 91.938 79.009 91.984 94.569 ;
        RECT 79.098 91.849 94.632 91.921 ;
        RECT 91.892 79.055 91.938 94.615 ;
        RECT 79.144 91.803 94.678 91.875 ;
        RECT 91.846 79.101 91.892 94.661 ;
        RECT 79.19 91.757 94.724 91.829 ;
        RECT 91.8 79.147 91.846 94.707 ;
        RECT 79.236 91.711 94.77 91.783 ;
        RECT 91.754 79.193 91.8 94.753 ;
        RECT 79.282 91.665 94.816 91.737 ;
        RECT 91.708 79.239 91.754 94.799 ;
        RECT 79.328 91.619 94.862 91.691 ;
        RECT 91.662 79.285 91.708 94.845 ;
        RECT 79.374 91.573 94.908 91.645 ;
        RECT 91.616 79.331 91.662 94.891 ;
        RECT 79.42 91.527 94.954 91.599 ;
        RECT 91.57 79.377 91.616 94.937 ;
        RECT 79.466 91.481 95 91.553 ;
        RECT 91.524 79.423 91.57 94.983 ;
        RECT 79.512 91.435 95.046 91.507 ;
        RECT 91.478 79.469 91.524 95.029 ;
        RECT 79.558 91.389 95.092 91.461 ;
        RECT 91.432 79.515 91.478 95.075 ;
        RECT 79.604 91.343 95.138 91.415 ;
        RECT 91.386 79.561 91.432 95.121 ;
        RECT 79.65 91.297 95.184 91.369 ;
        RECT 91.34 79.607 91.386 95.167 ;
        RECT 79.696 91.251 95.23 91.323 ;
        RECT 91.294 79.653 91.34 95.213 ;
        RECT 79.742 91.205 95.276 91.277 ;
        RECT 91.248 79.699 91.294 95.259 ;
        RECT 79.788 91.159 95.322 91.231 ;
        RECT 91.202 79.745 91.248 95.305 ;
        RECT 79.834 91.113 95.368 91.185 ;
        RECT 91.156 79.791 91.202 95.351 ;
        RECT 79.88 91.067 95.414 91.139 ;
        RECT 91.11 79.837 91.156 95.397 ;
        RECT 79.926 91.021 95.46 91.093 ;
        RECT 91.064 79.883 91.11 95.443 ;
        RECT 79.972 90.975 95.506 91.047 ;
        RECT 91.018 79.929 91.064 95.489 ;
        RECT 80.018 90.929 95.552 91.001 ;
        RECT 90.972 79.975 91.018 95.535 ;
        RECT 80.064 90.883 95.598 90.955 ;
        RECT 90.926 80.021 90.972 95.581 ;
        RECT 80.11 90.837 95.644 90.909 ;
        RECT 90.88 80.067 90.926 95.627 ;
        RECT 80.156 90.791 95.69 90.863 ;
        RECT 90.834 80.113 90.88 95.673 ;
        RECT 80.202 90.745 95.736 90.817 ;
        RECT 90.788 80.159 90.834 95.719 ;
        RECT 80.248 90.699 95.782 90.771 ;
        RECT 90.742 80.205 90.788 95.765 ;
        RECT 80.294 90.653 95.828 90.725 ;
        RECT 90.696 80.251 90.742 95.811 ;
        RECT 80.34 90.607 95.874 90.679 ;
        RECT 90.65 80.297 90.696 95.857 ;
        RECT 80.386 90.561 95.92 90.633 ;
        RECT 90.604 80.343 90.65 95.903 ;
        RECT 80.432 90.515 95.966 90.587 ;
        RECT 90.558 80.389 90.604 95.949 ;
        RECT 80.478 90.469 96.012 90.541 ;
        RECT 90.512 80.435 90.558 95.995 ;
        RECT 80.524 90.423 96.058 90.495 ;
        RECT 90.466 80.481 90.512 96.041 ;
        RECT 80.57 90.377 96.104 90.449 ;
        RECT 90.42 80.527 90.466 96.087 ;
        RECT 80.616 90.331 96.15 90.403 ;
        RECT 90.374 80.573 90.42 96.133 ;
        RECT 80.662 90.285 96.196 90.357 ;
        RECT 90.328 80.619 90.374 96.179 ;
        RECT 80.708 90.239 96.242 90.311 ;
        RECT 90.282 80.665 90.328 96.225 ;
        RECT 80.754 90.193 96.288 90.265 ;
        RECT 90.236 80.711 90.282 96.271 ;
        RECT 80.8 90.147 96.334 90.219 ;
        RECT 90.19 80.757 90.236 96.317 ;
        RECT 80.846 90.101 96.38 90.173 ;
        RECT 90.144 80.803 90.19 96.363 ;
        RECT 80.892 90.055 96.426 90.127 ;
        RECT 90.098 80.849 90.144 96.409 ;
        RECT 80.938 90.009 96.472 90.081 ;
        RECT 90.052 80.895 90.098 96.455 ;
        RECT 80.984 89.963 96.518 90.035 ;
        RECT 90.006 80.941 90.052 96.501 ;
        RECT 81.03 89.917 96.564 89.989 ;
        RECT 89.96 80.987 90.006 96.547 ;
        RECT 81.076 89.871 96.61 89.943 ;
        RECT 89.914 81.033 89.96 96.593 ;
        RECT 81.122 89.825 96.656 89.897 ;
        RECT 89.868 81.079 89.914 96.639 ;
        RECT 81.168 89.779 96.702 89.851 ;
        RECT 89.822 81.125 89.868 96.685 ;
        RECT 81.214 89.733 96.748 89.805 ;
        RECT 89.776 81.171 89.822 96.731 ;
        RECT 81.26 89.687 96.794 89.759 ;
        RECT 89.73 81.217 89.776 96.777 ;
        RECT 81.306 89.641 96.84 89.713 ;
        RECT 89.684 81.263 89.73 96.823 ;
        RECT 81.352 89.595 96.886 89.667 ;
        RECT 89.638 81.309 89.684 96.869 ;
        RECT 81.398 89.549 96.932 89.621 ;
        RECT 89.592 81.355 89.638 96.915 ;
        RECT 81.444 89.503 96.978 89.575 ;
        RECT 89.546 81.401 89.592 96.961 ;
        RECT 81.49 89.457 97.03 89.503 ;
        RECT 89.5 81.447 89.546 97.007 ;
        RECT 78.5 92.447 89.5 110 ;
        RECT 81.536 89.411 110 89.5 ;
        RECT 89.494 81.473 89.5 110 ;
        RECT 81.582 89.365 110 89.5 ;
        RECT 89.448 81.499 89.5 110 ;
        RECT 81.628 89.319 110 89.5 ;
        RECT 89.402 81.545 89.5 110 ;
        RECT 81.674 89.273 110 89.5 ;
        RECT 89.356 81.591 89.5 110 ;
        RECT 81.72 89.227 110 89.5 ;
        RECT 89.31 81.637 89.5 110 ;
        RECT 81.766 89.181 110 89.5 ;
        RECT 89.264 81.683 89.5 110 ;
        RECT 81.812 89.135 110 89.5 ;
        RECT 89.218 81.729 89.5 110 ;
        RECT 81.858 89.089 110 89.5 ;
        RECT 89.172 81.775 89.5 110 ;
        RECT 81.904 89.043 110 89.5 ;
        RECT 89.126 81.821 89.5 110 ;
        RECT 81.95 88.997 110 89.5 ;
        RECT 89.08 81.867 89.5 110 ;
        RECT 81.996 88.951 110 89.5 ;
        RECT 89.034 81.913 89.5 110 ;
        RECT 82.042 88.905 110 89.5 ;
        RECT 88.988 81.959 89.5 110 ;
        RECT 82.088 88.859 110 89.5 ;
        RECT 88.942 82.005 89.5 110 ;
        RECT 82.134 88.813 110 89.5 ;
        RECT 88.896 82.051 89.5 110 ;
        RECT 82.18 88.767 110 89.5 ;
        RECT 88.85 82.097 89.5 110 ;
        RECT 82.226 88.721 110 89.5 ;
        RECT 88.804 82.143 89.5 110 ;
        RECT 82.272 88.675 110 89.5 ;
        RECT 88.758 82.189 89.5 110 ;
        RECT 82.318 88.629 110 89.5 ;
        RECT 88.712 82.235 89.5 110 ;
        RECT 82.364 88.583 110 89.5 ;
        RECT 88.666 82.281 89.5 110 ;
        RECT 82.41 88.537 110 89.5 ;
        RECT 88.62 82.327 89.5 110 ;
        RECT 82.456 88.491 110 89.5 ;
        RECT 88.574 82.373 89.5 110 ;
        RECT 82.502 88.445 110 89.5 ;
        RECT 88.528 82.419 89.5 110 ;
        RECT 82.548 88.399 110 89.5 ;
        RECT 88.482 82.465 89.5 110 ;
        RECT 82.594 88.353 110 89.5 ;
        RECT 88.436 82.511 89.5 110 ;
        RECT 82.64 88.307 110 89.5 ;
        RECT 88.39 82.557 89.5 110 ;
        RECT 82.686 88.261 110 89.5 ;
        RECT 88.344 82.603 89.5 110 ;
        RECT 82.732 88.215 110 89.5 ;
        RECT 88.298 82.649 89.5 110 ;
        RECT 82.778 88.169 110 89.5 ;
        RECT 88.252 82.695 89.5 110 ;
        RECT 82.824 88.123 110 89.5 ;
        RECT 88.206 82.741 89.5 110 ;
        RECT 82.87 88.077 110 89.5 ;
        RECT 88.16 82.787 89.5 110 ;
        RECT 82.916 88.031 110 89.5 ;
        RECT 88.114 82.833 89.5 110 ;
        RECT 82.962 87.985 110 89.5 ;
        RECT 88.068 82.879 89.5 110 ;
        RECT 83.008 87.939 110 89.5 ;
        RECT 88.022 82.925 89.5 110 ;
        RECT 83.054 87.893 110 89.5 ;
        RECT 87.976 82.971 89.5 110 ;
        RECT 83.1 87.847 110 89.5 ;
        RECT 87.93 83.017 89.5 110 ;
        RECT 83.146 87.801 110 89.5 ;
        RECT 87.884 83.063 89.5 110 ;
        RECT 83.192 87.755 110 89.5 ;
        RECT 87.838 83.109 89.5 110 ;
        RECT 83.238 87.709 110 89.5 ;
        RECT 87.792 83.155 89.5 110 ;
        RECT 83.284 87.663 110 89.5 ;
        RECT 87.746 83.201 89.5 110 ;
        RECT 83.33 87.617 110 89.5 ;
        RECT 87.7 83.247 89.5 110 ;
        RECT 83.376 87.571 110 89.5 ;
        RECT 87.654 83.293 89.5 110 ;
        RECT 83.422 87.525 110 89.5 ;
        RECT 87.608 83.339 89.5 110 ;
        RECT 83.468 87.479 110 89.5 ;
        RECT 87.562 83.385 89.5 110 ;
        RECT 83.514 87.433 110 89.5 ;
        RECT 87.516 83.431 89.5 110 ;
        RECT 83.56 87.387 110 89.5 ;
        RECT 87.47 83.477 89.5 110 ;
        RECT 83.606 87.341 110 89.5 ;
        RECT 87.424 83.523 89.5 110 ;
        RECT 83.652 87.295 110 89.5 ;
        RECT 87.378 83.569 89.5 110 ;
        RECT 83.698 87.249 110 89.5 ;
        RECT 87.332 83.615 89.5 110 ;
        RECT 83.744 87.203 110 89.5 ;
        RECT 87.286 83.661 89.5 110 ;
        RECT 83.79 87.157 110 89.5 ;
        RECT 87.24 83.707 89.5 110 ;
        RECT 83.836 87.111 110 89.5 ;
        RECT 87.194 83.753 89.5 110 ;
        RECT 83.882 87.065 110 89.5 ;
        RECT 87.148 83.799 89.5 110 ;
        RECT 83.928 87.019 110 89.5 ;
        RECT 87.102 83.845 89.5 110 ;
        RECT 83.974 86.973 110 89.5 ;
        RECT 87.056 83.891 89.5 110 ;
        RECT 84.02 86.927 110 89.5 ;
        RECT 87.01 83.937 89.5 110 ;
        RECT 84.066 86.881 110 89.5 ;
        RECT 86.964 83.983 89.5 110 ;
        RECT 84.112 86.835 110 89.5 ;
        RECT 86.918 84.029 89.5 110 ;
        RECT 84.158 86.789 110 89.5 ;
        RECT 86.872 84.075 89.5 110 ;
        RECT 84.204 86.743 110 89.5 ;
        RECT 86.826 84.121 89.5 110 ;
        RECT 84.25 86.697 110 89.5 ;
        RECT 86.78 84.167 89.5 110 ;
        RECT 84.296 86.651 110 89.5 ;
        RECT 86.734 84.213 89.5 110 ;
        RECT 84.342 86.605 110 89.5 ;
        RECT 86.688 84.259 89.5 110 ;
        RECT 84.388 86.559 110 89.5 ;
        RECT 86.642 84.305 89.5 110 ;
        RECT 84.434 86.513 110 89.5 ;
        RECT 86.596 84.351 89.5 110 ;
        RECT 84.48 86.467 110 89.5 ;
        RECT 86.55 84.397 89.5 110 ;
        RECT 84.526 86.421 110 89.5 ;
        RECT 86.504 84.443 89.5 110 ;
        RECT 84.572 86.375 110 89.5 ;
        RECT 86.458 84.489 89.5 110 ;
        RECT 84.618 86.329 110 89.5 ;
        RECT 86.412 84.535 89.5 110 ;
        RECT 84.664 86.283 110 89.5 ;
        RECT 86.366 84.581 89.5 110 ;
        RECT 84.71 86.237 110 89.5 ;
        RECT 86.32 84.627 89.5 110 ;
        RECT 84.756 86.191 110 89.5 ;
        RECT 86.274 84.673 89.5 110 ;
        RECT 84.802 86.145 110 89.5 ;
        RECT 86.228 84.719 89.5 110 ;
        RECT 84.848 86.099 110 89.5 ;
        RECT 86.182 84.765 89.5 110 ;
        RECT 84.894 86.053 110 89.5 ;
        RECT 86.136 84.811 89.5 110 ;
        RECT 84.94 86.007 110 89.5 ;
        RECT 86.09 84.857 89.5 110 ;
        RECT 84.986 85.961 110 89.5 ;
        RECT 86.044 84.903 89.5 110 ;
        RECT 85.032 85.915 110 89.5 ;
        RECT 85.998 84.949 89.5 110 ;
        RECT 85.078 85.869 110 89.5 ;
        RECT 85.952 84.995 89.5 110 ;
        RECT 85.124 85.823 110 89.5 ;
        RECT 85.906 85.041 89.5 110 ;
        RECT 85.17 85.777 110 89.5 ;
        RECT 85.86 85.087 89.5 110 ;
        RECT 85.216 85.731 110 89.5 ;
        RECT 85.814 85.133 89.5 110 ;
        RECT 85.262 85.685 110 89.5 ;
        RECT 85.768 85.179 89.5 110 ;
        RECT 85.308 85.639 110 89.5 ;
        RECT 85.722 85.225 89.5 110 ;
        RECT 85.354 85.593 110 89.5 ;
        RECT 85.676 85.271 89.5 110 ;
        RECT 85.4 85.547 110 89.5 ;
        RECT 85.63 85.317 89.5 110 ;
        RECT 85.446 85.501 110 89.5 ;
        RECT 85.584 85.363 89.5 110 ;
        RECT 85.492 85.455 110 89.5 ;
        RECT 85.538 85.409 89.5 110 ;
        RECT 10.032 49.46 27 49.508 ;
        RECT 9.986 49.506 26.954 49.554 ;
        RECT 9.94 49.552 26.908 49.6 ;
        RECT 9.894 49.598 26.862 49.646 ;
        RECT 9.848 49.644 26.816 49.692 ;
        RECT 9.802 49.69 26.77 49.738 ;
        RECT 9.756 49.736 26.724 49.784 ;
        RECT 9.71 49.782 26.678 49.83 ;
        RECT 9.664 49.828 26.632 49.876 ;
        RECT 9.618 49.874 26.586 49.922 ;
        RECT 9.572 49.92 26.54 49.968 ;
        RECT 9.526 49.966 26.494 50.014 ;
        RECT 9.48 50.012 26.448 50.06 ;
        RECT 9.434 50.058 26.402 50.106 ;
        RECT 9.388 50.104 26.356 50.152 ;
        RECT 9.342 50.15 26.31 50.198 ;
        RECT 9.296 50.196 26.264 50.244 ;
        RECT 9.25 50.242 26.218 50.29 ;
        RECT 9.204 50.288 26.172 50.336 ;
        RECT 9.158 50.334 26.126 50.382 ;
        RECT 9.112 50.38 26.08 50.428 ;
        RECT 9.066 50.426 26.034 50.474 ;
        RECT 9.02 50.472 25.988 50.52 ;
        RECT 8.974 50.518 25.942 50.566 ;
        RECT 8.928 50.564 25.896 50.612 ;
        RECT 8.882 50.61 25.85 50.658 ;
        RECT 8.836 50.656 25.804 50.704 ;
        RECT 8.79 50.702 25.758 50.75 ;
        RECT 8.744 50.748 25.712 50.796 ;
        RECT 8.698 50.794 25.666 50.842 ;
        RECT 8.652 50.84 25.62 50.888 ;
        RECT 8.606 50.886 25.574 50.934 ;
        RECT 8.56 50.932 25.528 50.98 ;
        RECT 8.514 50.978 25.482 51.026 ;
        RECT 8.468 51.024 25.436 51.072 ;
        RECT 8.422 51.07 25.39 51.118 ;
        RECT 8.376 51.116 25.344 51.164 ;
        RECT 8.33 51.162 25.298 51.21 ;
        RECT 8.284 51.208 25.252 51.256 ;
        RECT 8.238 51.254 25.206 51.302 ;
        RECT 8.192 51.3 25.16 51.348 ;
        RECT 8.146 51.346 25.114 51.394 ;
        RECT 8.1 51.392 25.068 51.44 ;
        RECT 8.054 51.438 25.022 51.486 ;
        RECT 8.008 51.484 24.976 51.532 ;
        RECT 7.962 51.53 24.93 51.578 ;
        RECT 7.916 51.576 24.884 51.624 ;
        RECT 7.87 51.622 24.838 51.67 ;
        RECT 7.824 51.668 24.792 51.716 ;
        RECT 7.778 51.714 24.746 51.762 ;
        RECT 7.732 51.76 24.7 51.808 ;
        RECT 7.686 51.806 24.654 51.854 ;
        RECT 7.64 51.852 24.608 51.9 ;
        RECT 7.594 51.898 24.562 51.946 ;
        RECT 7.548 51.944 24.516 51.992 ;
        RECT 7.502 51.99 24.47 52.038 ;
        RECT 7.456 52.036 24.424 52.084 ;
        RECT 7.41 52.082 24.378 52.13 ;
        RECT 7.364 52.128 24.332 52.176 ;
        RECT 7.318 52.174 24.286 52.222 ;
        RECT 7.272 52.22 24.24 52.268 ;
        RECT 7.226 52.266 24.194 52.314 ;
        RECT 7.18 52.312 24.148 52.36 ;
        RECT 7.134 52.358 24.102 52.406 ;
        RECT 7.088 52.404 24.056 52.452 ;
        RECT 7.042 52.45 24.01 52.498 ;
        RECT 6.996 52.496 23.964 52.544 ;
        RECT 6.95 52.542 23.918 52.59 ;
        RECT 6.904 52.588 23.872 52.636 ;
        RECT 6.858 52.634 23.826 52.682 ;
        RECT 6.812 52.68 23.78 52.728 ;
        RECT 6.766 52.726 23.734 52.774 ;
        RECT 6.72 52.772 23.688 52.82 ;
        RECT 6.674 52.818 23.642 52.866 ;
        RECT 6.628 52.864 23.596 52.912 ;
        RECT 6.582 52.91 23.55 52.958 ;
        RECT 6.536 52.956 23.504 53.004 ;
        RECT 6.49 53.002 23.458 53.05 ;
        RECT 6.444 53.048 23.412 53.096 ;
        RECT 6.398 53.094 23.366 53.142 ;
        RECT 6.352 53.14 23.32 53.188 ;
        RECT 6.306 53.186 23.274 53.234 ;
        RECT 6.26 53.232 23.228 53.28 ;
        RECT 6.214 53.278 23.182 53.326 ;
        RECT 6.168 53.324 23.136 53.372 ;
        RECT 6.122 53.37 23.09 53.418 ;
        RECT 6.076 53.416 23.044 53.464 ;
        RECT 6.03 53.462 22.998 53.51 ;
        RECT 5.984 53.508 22.952 53.556 ;
        RECT 5.938 53.554 22.906 53.602 ;
        RECT 5.892 53.6 22.86 53.648 ;
        RECT 5.846 53.646 22.814 53.694 ;
        RECT 5.8 53.692 22.768 53.74 ;
        RECT 5.754 53.738 22.722 53.786 ;
        RECT 5.708 53.784 22.676 53.832 ;
        RECT 5.662 53.83 22.63 53.878 ;
        RECT 5.616 53.876 22.584 53.924 ;
        RECT 5.57 53.922 22.538 53.97 ;
        RECT 5.524 53.968 22.492 54.016 ;
        RECT 5.478 54.014 22.446 54.062 ;
        RECT 5.432 54.06 22.4 54.108 ;
        RECT 5.386 54.106 22.354 54.154 ;
        RECT 5.34 54.152 22.308 54.2 ;
        RECT 5.294 54.198 22.262 54.246 ;
        RECT 5.248 54.244 22.216 54.292 ;
        RECT 5.202 54.29 22.17 54.338 ;
        RECT 5.156 54.336 22.124 54.384 ;
        RECT 5.11 54.382 22.078 54.43 ;
        RECT 5.064 54.428 22.032 54.476 ;
        RECT 5.018 54.474 21.986 54.522 ;
        RECT 4.972 54.52 21.94 54.568 ;
        RECT 4.926 54.566 21.894 54.614 ;
        RECT 4.88 54.612 21.848 54.66 ;
        RECT 4.834 54.658 21.802 54.706 ;
        RECT 4.788 54.704 21.756 54.752 ;
        RECT 4.742 54.75 21.71 54.798 ;
        RECT 4.696 54.796 21.664 54.844 ;
        RECT 4.65 54.842 21.618 54.89 ;
        RECT 4.604 54.888 21.572 54.936 ;
        RECT 4.558 54.934 21.526 54.982 ;
        RECT 4.512 54.98 21.48 55.028 ;
        RECT 4.466 55.026 21.434 55.074 ;
        RECT 4.42 55.072 21.388 55.12 ;
        RECT 4.374 55.118 21.342 55.166 ;
        RECT 4.328 55.164 21.296 55.212 ;
        RECT 4.282 55.21 21.25 55.258 ;
        RECT 4.236 55.256 21.204 55.304 ;
        RECT 4.19 55.302 21.158 55.35 ;
        RECT 4.144 55.348 21.112 55.396 ;
        RECT 4.098 55.394 21.066 55.442 ;
        RECT 4.052 55.44 21.02 55.488 ;
        RECT 4.006 55.486 20.974 55.534 ;
        RECT 3.96 55.532 20.928 55.58 ;
        RECT 3.914 55.578 20.882 55.626 ;
        RECT 3.868 55.624 20.836 55.672 ;
        RECT 3.822 55.67 20.79 55.718 ;
        RECT 3.776 55.716 20.744 55.764 ;
        RECT 3.73 55.762 20.698 55.81 ;
        RECT 3.684 55.808 20.652 55.856 ;
        RECT 3.638 55.854 20.606 55.902 ;
        RECT 3.592 55.9 20.56 55.948 ;
        RECT 3.546 55.946 20.514 55.994 ;
        RECT 3.5 55.992 20.468 56.04 ;
        RECT 3.5 55.992 20.422 56.086 ;
        RECT 3.5 55.992 20.376 56.132 ;
        RECT 3.5 55.992 20.33 56.178 ;
        RECT 3.5 55.992 20.284 56.224 ;
        RECT 3.5 55.992 20.238 56.27 ;
        RECT 3.5 55.992 20.192 56.316 ;
        RECT 3.5 55.992 20.146 56.362 ;
        RECT 3.5 55.992 20.1 56.408 ;
        RECT 3.5 55.992 20.054 56.454 ;
        RECT 3.5 55.992 20.008 56.5 ;
        RECT 3.5 55.992 19.962 56.546 ;
        RECT 3.5 55.992 19.916 56.592 ;
        RECT 3.5 55.992 19.87 56.638 ;
        RECT 3.5 55.992 19.824 56.684 ;
        RECT 3.5 55.992 19.778 56.73 ;
        RECT 3.5 55.992 19.732 56.776 ;
        RECT 3.5 55.992 19.686 56.822 ;
        RECT 3.5 55.992 19.64 56.868 ;
        RECT 3.5 55.992 19.594 56.914 ;
        RECT 3.5 55.992 19.548 56.96 ;
        RECT 3.5 55.992 19.502 57.006 ;
        RECT 3.5 55.992 19.456 57.052 ;
        RECT 3.5 55.992 19.41 57.098 ;
        RECT 3.5 55.992 19.364 57.144 ;
        RECT 3.5 55.992 19.318 57.19 ;
        RECT 3.5 55.992 19.272 57.236 ;
        RECT 3.5 55.992 19.226 57.282 ;
        RECT 3.5 55.992 19.18 57.328 ;
        RECT 3.5 55.992 19.134 57.374 ;
        RECT 3.5 55.992 19.088 57.42 ;
        RECT 3.5 55.992 19.042 57.466 ;
        RECT 3.5 55.992 18.996 57.512 ;
        RECT 3.5 55.992 18.95 57.558 ;
        RECT 3.5 55.992 18.904 57.604 ;
        RECT 3.5 55.992 18.858 57.65 ;
        RECT 3.5 55.992 18.812 57.696 ;
        RECT 3.5 55.992 18.766 57.742 ;
        RECT 3.5 55.992 18.72 57.788 ;
        RECT 3.5 55.992 18.674 57.834 ;
        RECT 3.5 55.992 18.628 57.88 ;
        RECT 3.5 55.992 18.582 57.926 ;
        RECT 3.5 55.992 18.536 57.972 ;
        RECT 3.5 55.992 18.49 58.018 ;
        RECT 3.5 55.992 18.444 58.064 ;
        RECT 3.5 55.992 18.398 58.11 ;
        RECT 3.5 55.992 18.352 58.156 ;
        RECT 3.5 55.992 18.306 58.202 ;
        RECT 3.5 55.992 18.26 58.248 ;
        RECT 3.5 55.992 18.214 58.294 ;
        RECT 3.5 55.992 18.168 58.34 ;
        RECT 3.5 55.992 18.122 58.386 ;
        RECT 3.5 55.992 18.076 58.432 ;
        RECT 3.5 55.992 18.03 58.478 ;
        RECT 3.5 55.992 17.984 58.524 ;
        RECT 3.5 55.992 17.938 58.57 ;
        RECT 3.5 55.992 17.892 58.616 ;
        RECT 3.5 55.992 17.846 58.662 ;
        RECT 3.5 55.992 17.8 58.708 ;
        RECT 3.5 55.992 17.754 58.754 ;
        RECT 3.5 55.992 17.708 58.8 ;
        RECT 3.5 55.992 17.662 58.846 ;
        RECT 3.5 55.992 17.616 58.892 ;
        RECT 3.5 55.992 17.57 58.938 ;
        RECT 3.5 55.992 17.524 58.984 ;
        RECT 3.5 55.992 17.478 59.03 ;
        RECT 3.5 55.992 17.432 59.076 ;
        RECT 3.5 55.992 17.386 59.122 ;
        RECT 3.5 55.992 17.34 59.168 ;
        RECT 3.5 55.992 17.294 59.214 ;
        RECT 3.5 55.992 17.248 59.26 ;
        RECT 3.5 55.992 17.202 59.306 ;
        RECT 3.5 55.992 17.156 59.352 ;
        RECT 3.5 55.992 17.11 59.398 ;
        RECT 3.5 55.992 17.064 59.444 ;
        RECT 3.5 55.992 17.018 59.49 ;
        RECT 3.5 55.992 16.972 59.536 ;
        RECT 3.5 55.992 16.926 59.582 ;
        RECT 3.5 55.992 16.88 59.628 ;
        RECT 3.5 55.992 16.834 59.674 ;
        RECT 3.5 55.992 16.788 59.72 ;
        RECT 3.5 55.992 16.742 59.766 ;
        RECT 3.5 55.992 16.696 59.812 ;
        RECT 3.5 55.992 16.65 59.858 ;
        RECT 3.5 55.992 16.604 59.904 ;
        RECT 3.5 55.992 16.558 59.95 ;
        RECT 3.5 55.992 16.512 59.996 ;
        RECT 3.5 55.992 16.466 60.042 ;
        RECT 3.5 55.992 16.42 60.088 ;
        RECT 3.5 55.992 16.374 60.134 ;
        RECT 3.5 55.992 16.328 60.18 ;
        RECT 3.5 55.992 16.282 60.226 ;
        RECT 3.5 55.992 16.236 60.272 ;
        RECT 3.5 55.992 16.19 60.318 ;
        RECT 3.5 55.992 16.144 60.364 ;
        RECT 3.5 55.992 16.098 60.41 ;
        RECT 3.5 55.992 16.052 60.456 ;
        RECT 3.5 55.992 16.006 60.502 ;
        RECT 3.5 55.992 15.96 60.548 ;
        RECT 3.5 55.992 15.914 60.594 ;
        RECT 3.5 55.992 15.868 60.64 ;
        RECT 3.5 55.992 15.822 60.686 ;
        RECT 3.5 55.992 15.776 60.732 ;
        RECT 3.5 55.992 15.73 60.778 ;
        RECT 3.5 55.992 15.684 60.824 ;
        RECT 3.5 55.992 15.638 60.87 ;
        RECT 3.5 55.992 15.592 60.916 ;
        RECT 3.5 55.992 15.546 60.962 ;
        RECT 3.5 55.992 15.5 110 ;
        RECT 62.764 17 110 29 ;
        RECT 50.758 28.984 67.733 29.024 ;
        RECT 45.836 33.906 62.765 33.971 ;
        RECT 62.718 17.024 62.764 33.994 ;
        RECT 45.79 33.952 62.718 34.04 ;
        RECT 45.882 33.86 62.811 33.947 ;
        RECT 62.672 17.07 62.718 34.04 ;
        RECT 45.744 33.998 62.672 34.086 ;
        RECT 45.928 33.814 62.857 33.901 ;
        RECT 62.626 17.116 62.672 34.086 ;
        RECT 45.698 34.044 62.626 34.132 ;
        RECT 45.974 33.768 62.903 33.855 ;
        RECT 62.58 17.162 62.626 34.132 ;
        RECT 45.652 34.09 62.58 34.178 ;
        RECT 46.02 33.722 62.949 33.809 ;
        RECT 62.534 17.208 62.58 34.178 ;
        RECT 45.606 34.136 62.534 34.224 ;
        RECT 46.066 33.676 62.995 33.763 ;
        RECT 62.488 17.254 62.534 34.224 ;
        RECT 45.56 34.182 62.488 34.27 ;
        RECT 46.112 33.63 63.041 33.717 ;
        RECT 62.442 17.3 62.488 34.27 ;
        RECT 45.514 34.228 62.442 34.316 ;
        RECT 46.158 33.584 63.087 33.671 ;
        RECT 62.396 17.346 62.442 34.316 ;
        RECT 45.468 34.274 62.396 34.362 ;
        RECT 46.204 33.538 63.133 33.625 ;
        RECT 62.35 17.392 62.396 34.362 ;
        RECT 45.422 34.32 62.35 34.408 ;
        RECT 46.25 33.492 63.179 33.579 ;
        RECT 62.304 17.438 62.35 34.408 ;
        RECT 45.376 34.366 62.304 34.454 ;
        RECT 46.296 33.446 63.225 33.533 ;
        RECT 62.258 17.484 62.304 34.454 ;
        RECT 45.33 34.412 62.258 34.5 ;
        RECT 46.342 33.4 63.271 33.487 ;
        RECT 62.212 17.53 62.258 34.5 ;
        RECT 45.284 34.458 62.212 34.546 ;
        RECT 46.388 33.354 63.317 33.441 ;
        RECT 62.166 17.576 62.212 34.546 ;
        RECT 45.238 34.504 62.166 34.592 ;
        RECT 46.434 33.308 63.363 33.395 ;
        RECT 62.12 17.622 62.166 34.592 ;
        RECT 45.192 34.55 62.12 34.638 ;
        RECT 46.48 33.262 63.409 33.349 ;
        RECT 62.074 17.668 62.12 34.638 ;
        RECT 45.146 34.596 62.074 34.684 ;
        RECT 46.526 33.216 63.455 33.303 ;
        RECT 62.028 17.714 62.074 34.684 ;
        RECT 45.1 34.642 62.028 34.73 ;
        RECT 46.572 33.17 63.501 33.257 ;
        RECT 61.982 17.76 62.028 34.73 ;
        RECT 45.054 34.688 61.982 34.776 ;
        RECT 46.618 33.124 63.547 33.211 ;
        RECT 61.936 17.806 61.982 34.776 ;
        RECT 45.008 34.734 61.936 34.822 ;
        RECT 46.664 33.078 63.593 33.165 ;
        RECT 61.89 17.852 61.936 34.822 ;
        RECT 44.962 34.78 61.89 34.868 ;
        RECT 46.71 33.032 63.639 33.119 ;
        RECT 61.844 17.898 61.89 34.868 ;
        RECT 44.916 34.826 61.844 34.914 ;
        RECT 46.756 32.986 63.685 33.073 ;
        RECT 61.798 17.944 61.844 34.914 ;
        RECT 44.87 34.872 61.798 34.96 ;
        RECT 46.802 32.94 63.731 33.027 ;
        RECT 61.752 17.99 61.798 34.96 ;
        RECT 44.824 34.918 61.752 35.006 ;
        RECT 46.848 32.894 63.777 32.981 ;
        RECT 61.706 18.036 61.752 35.006 ;
        RECT 44.778 34.964 61.706 35.052 ;
        RECT 46.894 32.848 63.823 32.935 ;
        RECT 61.66 18.082 61.706 35.052 ;
        RECT 44.732 35.01 61.66 35.098 ;
        RECT 46.94 32.802 63.869 32.889 ;
        RECT 61.614 18.128 61.66 35.098 ;
        RECT 44.686 35.056 61.614 35.144 ;
        RECT 46.986 32.756 63.915 32.843 ;
        RECT 61.568 18.174 61.614 35.144 ;
        RECT 44.64 35.102 61.568 35.19 ;
        RECT 47.032 32.71 63.961 32.797 ;
        RECT 61.522 18.22 61.568 35.19 ;
        RECT 44.594 35.148 61.522 35.236 ;
        RECT 47.078 32.664 64.007 32.751 ;
        RECT 61.476 18.266 61.522 35.236 ;
        RECT 44.548 35.194 61.476 35.282 ;
        RECT 47.124 32.618 64.053 32.705 ;
        RECT 61.43 18.312 61.476 35.282 ;
        RECT 44.502 35.24 61.43 35.328 ;
        RECT 47.17 32.572 64.099 32.659 ;
        RECT 61.384 18.358 61.43 35.328 ;
        RECT 44.456 35.286 61.384 35.374 ;
        RECT 47.216 32.526 64.145 32.613 ;
        RECT 61.338 18.404 61.384 35.374 ;
        RECT 44.41 35.332 61.338 35.42 ;
        RECT 47.262 32.48 64.191 32.567 ;
        RECT 61.292 18.45 61.338 35.42 ;
        RECT 44.364 35.378 61.292 35.466 ;
        RECT 47.308 32.434 64.237 32.521 ;
        RECT 61.246 18.496 61.292 35.466 ;
        RECT 44.318 35.424 61.246 35.512 ;
        RECT 47.354 32.388 64.283 32.475 ;
        RECT 61.2 18.542 61.246 35.512 ;
        RECT 44.272 35.47 61.2 35.558 ;
        RECT 47.4 32.342 64.329 32.429 ;
        RECT 61.154 18.588 61.2 35.558 ;
        RECT 44.226 35.516 61.154 35.604 ;
        RECT 47.446 32.296 64.375 32.383 ;
        RECT 61.108 18.634 61.154 35.604 ;
        RECT 44.18 35.562 61.108 35.65 ;
        RECT 47.492 32.25 64.421 32.337 ;
        RECT 61.062 18.68 61.108 35.65 ;
        RECT 44.134 35.608 61.062 35.696 ;
        RECT 47.538 32.204 64.467 32.291 ;
        RECT 61.016 18.726 61.062 35.696 ;
        RECT 44.088 35.654 61.016 35.742 ;
        RECT 47.584 32.158 64.513 32.245 ;
        RECT 60.97 18.772 61.016 35.742 ;
        RECT 44.042 35.7 60.97 35.788 ;
        RECT 47.63 32.112 64.559 32.199 ;
        RECT 60.924 18.818 60.97 35.788 ;
        RECT 43.996 35.746 60.924 35.834 ;
        RECT 47.676 32.066 64.605 32.153 ;
        RECT 60.878 18.864 60.924 35.834 ;
        RECT 43.95 35.792 60.878 35.88 ;
        RECT 47.722 32.02 64.651 32.107 ;
        RECT 60.832 18.91 60.878 35.88 ;
        RECT 43.904 35.838 60.832 35.926 ;
        RECT 47.768 31.974 64.697 32.061 ;
        RECT 60.786 18.956 60.832 35.926 ;
        RECT 43.858 35.884 60.786 35.972 ;
        RECT 47.814 31.928 64.743 32.015 ;
        RECT 60.74 19.002 60.786 35.972 ;
        RECT 43.812 35.93 60.74 36.018 ;
        RECT 47.86 31.882 64.789 31.969 ;
        RECT 60.694 19.048 60.74 36.018 ;
        RECT 43.766 35.976 60.694 36.064 ;
        RECT 47.906 31.836 64.835 31.923 ;
        RECT 60.648 19.094 60.694 36.064 ;
        RECT 43.72 36.022 60.648 36.11 ;
        RECT 47.952 31.79 64.881 31.877 ;
        RECT 60.602 19.14 60.648 36.11 ;
        RECT 43.674 36.068 60.602 36.156 ;
        RECT 47.998 31.744 64.927 31.831 ;
        RECT 60.556 19.186 60.602 36.156 ;
        RECT 43.628 36.114 60.556 36.202 ;
        RECT 48.044 31.698 64.973 31.785 ;
        RECT 60.51 19.232 60.556 36.202 ;
        RECT 43.582 36.16 60.51 36.248 ;
        RECT 48.09 31.652 65.019 31.739 ;
        RECT 60.464 19.278 60.51 36.248 ;
        RECT 43.536 36.206 60.464 36.294 ;
        RECT 48.136 31.606 65.065 31.693 ;
        RECT 60.418 19.324 60.464 36.294 ;
        RECT 43.49 36.252 60.418 36.34 ;
        RECT 48.182 31.56 65.111 31.647 ;
        RECT 60.372 19.37 60.418 36.34 ;
        RECT 43.444 36.298 60.372 36.386 ;
        RECT 48.228 31.514 65.157 31.601 ;
        RECT 60.326 19.416 60.372 36.386 ;
        RECT 43.398 36.344 60.326 36.432 ;
        RECT 48.274 31.468 65.203 31.555 ;
        RECT 60.28 19.462 60.326 36.432 ;
        RECT 43.352 36.39 60.28 36.478 ;
        RECT 48.32 31.422 65.249 31.509 ;
        RECT 60.234 19.508 60.28 36.478 ;
        RECT 43.306 36.436 60.234 36.524 ;
        RECT 48.366 31.376 65.295 31.463 ;
        RECT 60.188 19.554 60.234 36.524 ;
        RECT 43.26 36.482 60.188 36.57 ;
        RECT 48.412 31.33 65.341 31.417 ;
        RECT 60.142 19.6 60.188 36.57 ;
        RECT 43.214 36.528 60.142 36.616 ;
        RECT 48.458 31.284 65.387 31.371 ;
        RECT 60.096 19.646 60.142 36.616 ;
        RECT 43.168 36.574 60.096 36.662 ;
        RECT 48.504 31.238 65.433 31.325 ;
        RECT 60.05 19.692 60.096 36.662 ;
        RECT 43.122 36.62 60.05 36.708 ;
        RECT 48.55 31.192 65.479 31.279 ;
        RECT 60.004 19.738 60.05 36.708 ;
        RECT 43.076 36.666 60.004 36.754 ;
        RECT 48.596 31.146 65.525 31.233 ;
        RECT 59.958 19.784 60.004 36.754 ;
        RECT 43.03 36.712 59.958 36.8 ;
        RECT 48.642 31.1 65.571 31.187 ;
        RECT 59.912 19.83 59.958 36.8 ;
        RECT 42.984 36.758 59.912 36.846 ;
        RECT 48.688 31.054 65.617 31.141 ;
        RECT 59.866 19.876 59.912 36.846 ;
        RECT 42.938 36.804 59.866 36.892 ;
        RECT 48.734 31.008 65.663 31.095 ;
        RECT 59.82 19.922 59.866 36.892 ;
        RECT 42.892 36.85 59.82 36.938 ;
        RECT 48.78 30.962 65.709 31.049 ;
        RECT 59.774 19.968 59.82 36.938 ;
        RECT 42.846 36.896 59.774 36.984 ;
        RECT 48.826 30.916 65.755 31.003 ;
        RECT 59.728 20.014 59.774 36.984 ;
        RECT 42.8 36.942 59.728 37.03 ;
        RECT 48.872 30.87 65.801 30.957 ;
        RECT 59.682 20.06 59.728 37.03 ;
        RECT 42.754 36.988 59.682 37.076 ;
        RECT 48.918 30.824 65.847 30.911 ;
        RECT 59.636 20.106 59.682 37.076 ;
        RECT 42.708 37.034 59.636 37.122 ;
        RECT 48.964 30.778 65.893 30.865 ;
        RECT 59.59 20.152 59.636 37.122 ;
        RECT 42.662 37.08 59.59 37.168 ;
        RECT 49.01 30.732 65.939 30.819 ;
        RECT 59.544 20.198 59.59 37.168 ;
        RECT 42.616 37.126 59.544 37.214 ;
        RECT 49.056 30.686 65.985 30.773 ;
        RECT 59.498 20.244 59.544 37.214 ;
        RECT 42.57 37.172 59.498 37.26 ;
        RECT 49.102 30.64 66.031 30.727 ;
        RECT 59.452 20.29 59.498 37.26 ;
        RECT 42.524 37.218 59.452 37.306 ;
        RECT 49.148 30.594 66.077 30.681 ;
        RECT 59.406 20.336 59.452 37.306 ;
        RECT 42.478 37.264 59.406 37.352 ;
        RECT 49.194 30.548 66.123 30.635 ;
        RECT 59.36 20.382 59.406 37.352 ;
        RECT 42.432 37.31 59.36 37.398 ;
        RECT 49.24 30.502 66.169 30.589 ;
        RECT 59.314 20.428 59.36 37.398 ;
        RECT 42.386 37.356 59.314 37.444 ;
        RECT 49.286 30.456 66.215 30.543 ;
        RECT 59.268 20.474 59.314 37.444 ;
        RECT 42.34 37.402 59.268 37.49 ;
        RECT 49.332 30.41 66.261 30.497 ;
        RECT 59.222 20.52 59.268 37.49 ;
        RECT 42.294 37.448 59.222 37.536 ;
        RECT 49.378 30.364 66.307 30.451 ;
        RECT 59.176 20.566 59.222 37.536 ;
        RECT 42.248 37.494 59.176 37.582 ;
        RECT 49.424 30.318 66.353 30.405 ;
        RECT 59.13 20.612 59.176 37.582 ;
        RECT 42.202 37.54 59.13 37.628 ;
        RECT 49.47 30.272 66.399 30.359 ;
        RECT 59.084 20.658 59.13 37.628 ;
        RECT 42.156 37.586 59.084 37.674 ;
        RECT 49.516 30.226 66.445 30.313 ;
        RECT 59.038 20.704 59.084 37.674 ;
        RECT 42.11 37.632 59.038 37.72 ;
        RECT 49.562 30.18 66.491 30.267 ;
        RECT 58.992 20.75 59.038 37.72 ;
        RECT 42.064 37.678 58.992 37.766 ;
        RECT 49.608 30.134 66.537 30.221 ;
        RECT 58.946 20.796 58.992 37.766 ;
        RECT 42.018 37.724 58.946 37.812 ;
        RECT 49.654 30.088 66.583 30.175 ;
        RECT 58.9 20.842 58.946 37.812 ;
        RECT 41.972 37.77 58.9 37.858 ;
        RECT 49.7 30.042 66.629 30.129 ;
        RECT 58.854 20.888 58.9 37.858 ;
        RECT 41.926 37.816 58.854 37.904 ;
        RECT 49.746 29.996 66.675 30.083 ;
        RECT 58.808 20.934 58.854 37.904 ;
        RECT 41.88 37.862 58.808 37.95 ;
        RECT 49.792 29.95 66.721 30.037 ;
        RECT 58.762 20.98 58.808 37.95 ;
        RECT 41.834 37.908 58.762 37.996 ;
        RECT 49.838 29.904 66.767 29.991 ;
        RECT 58.716 21.026 58.762 37.996 ;
        RECT 41.788 37.954 58.716 38.042 ;
        RECT 49.884 29.858 66.813 29.945 ;
        RECT 58.67 21.072 58.716 38.042 ;
        RECT 41.742 38 58.67 38.088 ;
        RECT 49.93 29.812 66.859 29.899 ;
        RECT 58.624 21.118 58.67 38.088 ;
        RECT 41.696 38.046 58.624 38.134 ;
        RECT 49.976 29.766 66.905 29.853 ;
        RECT 58.578 21.164 58.624 38.134 ;
        RECT 41.65 38.092 58.578 38.18 ;
        RECT 50.022 29.72 66.951 29.807 ;
        RECT 58.532 21.21 58.578 38.18 ;
        RECT 41.604 38.138 58.532 38.226 ;
        RECT 50.068 29.674 66.997 29.761 ;
        RECT 58.486 21.256 58.532 38.226 ;
        RECT 41.558 38.184 58.486 38.272 ;
        RECT 50.114 29.628 67.043 29.715 ;
        RECT 58.44 21.302 58.486 38.272 ;
        RECT 41.512 38.23 58.44 38.318 ;
        RECT 50.16 29.582 67.089 29.669 ;
        RECT 58.394 21.348 58.44 38.318 ;
        RECT 41.466 38.276 58.394 38.364 ;
        RECT 50.206 29.536 67.135 29.623 ;
        RECT 58.348 21.394 58.394 38.364 ;
        RECT 41.42 38.322 58.348 38.41 ;
        RECT 50.252 29.49 67.181 29.577 ;
        RECT 58.302 21.44 58.348 38.41 ;
        RECT 41.374 38.368 58.302 38.456 ;
        RECT 50.298 29.444 67.227 29.531 ;
        RECT 58.256 21.486 58.302 38.456 ;
        RECT 41.328 38.414 58.256 38.502 ;
        RECT 50.344 29.398 67.273 29.485 ;
        RECT 58.21 21.532 58.256 38.502 ;
        RECT 41.282 38.46 58.21 38.548 ;
        RECT 50.39 29.352 67.319 29.439 ;
        RECT 58.164 21.578 58.21 38.548 ;
        RECT 41.236 38.506 58.164 38.594 ;
        RECT 50.436 29.306 67.365 29.393 ;
        RECT 58.118 21.624 58.164 38.594 ;
        RECT 41.19 38.552 58.118 38.64 ;
        RECT 50.482 29.26 67.411 29.347 ;
        RECT 58.072 21.67 58.118 38.64 ;
        RECT 41.144 38.598 58.072 38.686 ;
        RECT 50.528 29.214 67.457 29.301 ;
        RECT 58.026 21.716 58.072 38.686 ;
        RECT 41.098 38.644 58.026 38.732 ;
        RECT 50.574 29.168 67.503 29.255 ;
        RECT 57.98 21.762 58.026 38.732 ;
        RECT 41.052 38.69 57.98 38.778 ;
        RECT 50.62 29.122 67.549 29.209 ;
        RECT 57.934 21.808 57.98 38.778 ;
        RECT 41.006 38.736 57.934 38.824 ;
        RECT 50.666 29.076 67.595 29.163 ;
        RECT 57.888 21.854 57.934 38.824 ;
        RECT 40.96 38.782 57.888 38.87 ;
        RECT 50.712 29.03 67.641 29.117 ;
        RECT 57.842 21.9 57.888 38.87 ;
        RECT 40.914 38.828 57.842 38.916 ;
        RECT 50.758 28.984 67.687 29.071 ;
        RECT 57.796 21.946 57.842 38.916 ;
        RECT 40.868 38.874 57.796 38.962 ;
        RECT 50.804 28.938 110 29 ;
        RECT 57.75 21.992 57.796 38.962 ;
        RECT 40.822 38.92 57.75 39.008 ;
        RECT 50.85 28.892 110 29 ;
        RECT 57.704 22.038 57.75 39.008 ;
        RECT 40.776 38.966 57.704 39.054 ;
        RECT 50.896 28.846 110 29 ;
        RECT 57.658 22.084 57.704 39.054 ;
        RECT 40.73 39.012 57.658 39.1 ;
        RECT 50.942 28.8 110 29 ;
        RECT 57.612 22.13 57.658 39.1 ;
        RECT 40.684 39.058 57.612 39.146 ;
        RECT 50.988 28.754 110 29 ;
        RECT 57.566 22.176 57.612 39.146 ;
        RECT 40.638 39.104 57.566 39.192 ;
        RECT 51.034 28.708 110 29 ;
        RECT 57.52 22.222 57.566 39.192 ;
        RECT 40.592 39.15 57.52 39.238 ;
        RECT 51.08 28.662 110 29 ;
        RECT 57.474 22.268 57.52 39.238 ;
        RECT 40.546 39.196 57.474 39.284 ;
        RECT 51.126 28.616 110 29 ;
        RECT 57.428 22.314 57.474 39.284 ;
        RECT 40.5 39.242 57.428 39.33 ;
        RECT 51.172 28.57 110 29 ;
        RECT 57.382 22.36 57.428 39.33 ;
        RECT 40.454 39.288 57.382 39.376 ;
        RECT 51.218 28.524 110 29 ;
        RECT 57.336 22.406 57.382 39.376 ;
        RECT 40.408 39.334 57.336 39.422 ;
        RECT 51.264 28.478 110 29 ;
        RECT 57.29 22.452 57.336 39.422 ;
        RECT 40.362 39.38 57.29 39.468 ;
        RECT 51.31 28.432 110 29 ;
        RECT 57.244 22.498 57.29 39.468 ;
        RECT 40.316 39.426 57.244 39.514 ;
        RECT 51.356 28.386 110 29 ;
        RECT 57.198 22.544 57.244 39.514 ;
        RECT 40.27 39.472 57.198 39.56 ;
        RECT 51.402 28.34 110 29 ;
        RECT 57.152 22.59 57.198 39.56 ;
        RECT 40.224 39.518 57.152 39.606 ;
        RECT 51.448 28.294 110 29 ;
        RECT 57.106 22.636 57.152 39.606 ;
        RECT 40.178 39.564 57.106 39.652 ;
        RECT 51.494 28.248 110 29 ;
        RECT 57.06 22.682 57.106 39.652 ;
        RECT 40.132 39.61 57.06 39.698 ;
        RECT 51.54 28.202 110 29 ;
        RECT 57.014 22.728 57.06 39.698 ;
        RECT 40.086 39.656 57.014 39.744 ;
        RECT 51.586 28.156 110 29 ;
        RECT 56.968 22.774 57.014 39.744 ;
        RECT 40.04 39.702 56.968 39.79 ;
        RECT 51.632 28.11 110 29 ;
        RECT 56.922 22.82 56.968 39.79 ;
        RECT 39.994 39.748 56.922 39.836 ;
        RECT 51.678 28.064 110 29 ;
        RECT 56.876 22.866 56.922 39.836 ;
        RECT 39.948 39.794 56.876 39.882 ;
        RECT 51.724 28.018 110 29 ;
        RECT 56.83 22.912 56.876 39.882 ;
        RECT 39.902 39.84 56.83 39.928 ;
        RECT 51.77 27.972 110 29 ;
        RECT 56.784 22.958 56.83 39.928 ;
        RECT 39.856 39.886 56.784 39.974 ;
        RECT 51.816 27.926 110 29 ;
        RECT 56.738 23.004 56.784 39.974 ;
        RECT 39.81 39.932 56.738 40.02 ;
        RECT 51.862 27.88 110 29 ;
        RECT 56.692 23.05 56.738 40.02 ;
        RECT 39.764 39.978 56.692 40.066 ;
        RECT 51.908 27.834 110 29 ;
        RECT 56.646 23.096 56.692 40.066 ;
        RECT 39.718 40.024 56.646 40.112 ;
        RECT 51.954 27.788 110 29 ;
        RECT 56.6 23.142 56.646 40.112 ;
        RECT 39.672 40.07 56.6 40.158 ;
        RECT 52 27.742 110 29 ;
        RECT 56.554 23.188 56.6 40.158 ;
        RECT 39.626 40.116 56.554 40.204 ;
        RECT 52.046 27.696 110 29 ;
        RECT 56.508 23.234 56.554 40.204 ;
        RECT 39.58 40.162 56.508 40.25 ;
        RECT 52.092 27.65 110 29 ;
        RECT 56.462 23.28 56.508 40.25 ;
        RECT 39.534 40.208 56.462 40.296 ;
        RECT 52.138 27.604 110 29 ;
        RECT 56.416 23.326 56.462 40.296 ;
        RECT 39.488 40.254 56.416 40.342 ;
        RECT 52.184 27.558 110 29 ;
        RECT 56.37 23.372 56.416 40.342 ;
        RECT 39.442 40.3 56.37 40.388 ;
        RECT 52.23 27.512 110 29 ;
        RECT 56.324 23.418 56.37 40.388 ;
        RECT 39.396 40.346 56.324 40.434 ;
        RECT 52.276 27.466 110 29 ;
        RECT 56.278 23.464 56.324 40.434 ;
        RECT 39.35 40.392 56.278 40.48 ;
        RECT 52.322 27.42 110 29 ;
        RECT 56.232 23.51 56.278 40.48 ;
        RECT 39.304 40.438 56.232 40.526 ;
        RECT 52.368 27.374 110 29 ;
        RECT 56.186 23.556 56.232 40.526 ;
        RECT 39.258 40.484 56.186 40.572 ;
        RECT 52.414 27.328 110 29 ;
        RECT 56.14 23.602 56.186 40.572 ;
        RECT 39.212 40.53 56.14 40.618 ;
        RECT 52.46 27.282 110 29 ;
        RECT 56.094 23.648 56.14 40.618 ;
        RECT 39.166 40.576 56.094 40.664 ;
        RECT 52.506 27.236 110 29 ;
        RECT 56.048 23.694 56.094 40.664 ;
        RECT 39.12 40.622 56.048 40.71 ;
        RECT 52.552 27.19 110 29 ;
        RECT 56.002 23.74 56.048 40.71 ;
        RECT 39.074 40.668 56.002 40.756 ;
        RECT 52.598 27.144 110 29 ;
        RECT 55.956 23.786 56.002 40.756 ;
        RECT 39.028 40.714 55.956 40.802 ;
        RECT 52.644 27.098 110 29 ;
        RECT 55.91 23.832 55.956 40.802 ;
        RECT 38.982 40.76 55.91 40.848 ;
        RECT 52.69 27.052 110 29 ;
        RECT 55.864 23.878 55.91 40.848 ;
        RECT 38.936 40.806 55.864 40.894 ;
        RECT 52.736 27.006 110 29 ;
        RECT 55.818 23.924 55.864 40.894 ;
        RECT 38.89 40.852 55.818 40.94 ;
        RECT 52.782 26.96 110 29 ;
        RECT 55.772 23.97 55.818 40.94 ;
        RECT 38.844 40.898 55.772 40.986 ;
        RECT 52.828 26.914 110 29 ;
        RECT 55.726 24.016 55.772 40.986 ;
        RECT 38.798 40.944 55.726 41.032 ;
        RECT 52.874 26.868 110 29 ;
        RECT 55.68 24.062 55.726 41.032 ;
        RECT 38.752 40.99 55.68 41.078 ;
        RECT 52.92 26.822 110 29 ;
        RECT 55.634 24.108 55.68 41.078 ;
        RECT 38.706 41.036 55.634 41.124 ;
        RECT 52.966 26.776 110 29 ;
        RECT 55.588 24.154 55.634 41.124 ;
        RECT 38.66 41.082 55.588 41.17 ;
        RECT 53.012 26.73 110 29 ;
        RECT 55.542 24.2 55.588 41.17 ;
        RECT 38.614 41.128 55.542 41.216 ;
        RECT 53.058 26.684 110 29 ;
        RECT 55.496 24.246 55.542 41.216 ;
        RECT 38.568 41.174 55.496 41.262 ;
        RECT 53.104 26.638 110 29 ;
        RECT 55.45 24.292 55.496 41.262 ;
        RECT 38.522 41.22 55.45 41.308 ;
        RECT 53.15 26.592 110 29 ;
        RECT 55.404 24.338 55.45 41.308 ;
        RECT 38.476 41.266 55.404 41.354 ;
        RECT 53.196 26.546 110 29 ;
        RECT 55.358 24.384 55.404 41.354 ;
        RECT 38.43 41.312 55.358 41.4 ;
        RECT 53.242 26.5 110 29 ;
        RECT 55.312 24.43 55.358 41.4 ;
        RECT 38.384 41.358 55.312 41.446 ;
        RECT 53.288 26.454 110 29 ;
        RECT 55.266 24.476 55.312 41.446 ;
        RECT 38.338 41.404 55.266 41.492 ;
        RECT 53.334 26.408 110 29 ;
        RECT 55.22 24.522 55.266 41.492 ;
        RECT 38.292 41.45 55.22 41.538 ;
        RECT 53.38 26.362 110 29 ;
        RECT 55.174 24.568 55.22 41.538 ;
        RECT 38.246 41.496 55.174 41.584 ;
        RECT 53.426 26.316 110 29 ;
        RECT 55.128 24.614 55.174 41.584 ;
        RECT 38.2 41.542 55.128 41.63 ;
        RECT 53.472 26.27 110 29 ;
        RECT 55.082 24.66 55.128 41.63 ;
        RECT 38.154 41.588 55.082 41.676 ;
        RECT 53.518 26.224 110 29 ;
        RECT 55.036 24.706 55.082 41.676 ;
        RECT 38.108 41.634 55.036 41.722 ;
        RECT 53.564 26.178 110 29 ;
        RECT 54.99 24.752 55.036 41.722 ;
        RECT 38.062 41.68 54.99 41.768 ;
        RECT 53.61 26.132 110 29 ;
        RECT 54.944 24.798 54.99 41.768 ;
        RECT 38.016 41.726 54.944 41.814 ;
        RECT 53.656 26.086 110 29 ;
        RECT 54.898 24.844 54.944 41.814 ;
        RECT 37.97 41.772 54.898 41.86 ;
        RECT 53.702 26.04 110 29 ;
        RECT 54.852 24.89 54.898 41.86 ;
        RECT 37.924 41.818 54.852 41.906 ;
        RECT 53.748 25.994 110 29 ;
        RECT 54.806 24.936 54.852 41.906 ;
        RECT 37.878 41.864 54.806 41.952 ;
        RECT 53.794 25.948 110 29 ;
        RECT 54.76 24.982 54.806 41.952 ;
        RECT 37.832 41.91 54.76 41.998 ;
        RECT 53.84 25.902 110 29 ;
        RECT 54.714 25.028 54.76 41.998 ;
        RECT 37.786 41.956 54.714 42.044 ;
        RECT 53.886 25.856 110 29 ;
        RECT 54.668 25.074 54.714 42.044 ;
        RECT 37.74 42.002 54.668 42.09 ;
        RECT 53.932 25.81 110 29 ;
        RECT 54.622 25.12 54.668 42.09 ;
        RECT 37.694 42.048 54.622 42.136 ;
        RECT 53.978 25.764 110 29 ;
        RECT 54.576 25.166 54.622 42.136 ;
        RECT 37.648 42.094 54.576 42.182 ;
        RECT 54.024 25.718 110 29 ;
        RECT 54.53 25.212 54.576 42.182 ;
        RECT 37.602 42.14 54.53 42.228 ;
        RECT 54.07 25.672 110 29 ;
        RECT 54.484 25.258 54.53 42.228 ;
        RECT 37.556 42.186 54.484 42.274 ;
        RECT 54.116 25.626 110 29 ;
        RECT 54.438 25.304 54.484 42.274 ;
        RECT 37.51 42.232 54.438 42.32 ;
        RECT 54.162 25.58 110 29 ;
        RECT 54.392 25.35 54.438 42.32 ;
        RECT 37.464 42.278 54.392 42.366 ;
        RECT 54.208 25.534 110 29 ;
        RECT 54.346 25.396 54.392 42.366 ;
        RECT 37.418 42.324 54.346 42.412 ;
        RECT 54.254 25.488 110 29 ;
        RECT 54.3 25.442 54.346 42.412 ;
        RECT 37.372 42.37 54.3 42.458 ;
        RECT 37.326 42.416 54.254 42.504 ;
        RECT 37.28 42.462 54.208 42.55 ;
        RECT 37.234 42.508 54.162 42.596 ;
        RECT 37.188 42.554 54.116 42.642 ;
        RECT 37.142 42.6 54.07 42.688 ;
        RECT 37.096 42.646 54.024 42.734 ;
        RECT 37.05 42.692 53.978 42.78 ;
        RECT 37.004 42.738 53.932 42.826 ;
        RECT 36.958 42.784 53.886 42.872 ;
        RECT 36.912 42.83 53.84 42.918 ;
        RECT 36.866 42.876 53.794 42.964 ;
        RECT 36.82 42.922 53.748 43.01 ;
        RECT 36.774 42.968 53.702 43.056 ;
        RECT 36.728 43.014 53.656 43.102 ;
        RECT 36.682 43.06 53.61 43.148 ;
        RECT 36.636 43.106 53.564 43.194 ;
        RECT 36.59 43.152 53.518 43.24 ;
        RECT 36.544 43.198 53.472 43.286 ;
        RECT 36.498 43.244 53.426 43.332 ;
        RECT 36.452 43.29 53.38 43.378 ;
        RECT 36.406 43.336 53.334 43.424 ;
        RECT 36.36 43.382 53.288 43.47 ;
        RECT 36.314 43.428 53.242 43.516 ;
        RECT 36.268 43.474 53.196 43.562 ;
        RECT 36.222 43.52 53.15 43.608 ;
        RECT 36.176 43.566 53.104 43.654 ;
        RECT 36.13 43.612 53.058 43.7 ;
        RECT 36.084 43.658 53.012 43.746 ;
        RECT 36.038 43.704 52.966 43.792 ;
        RECT 35.992 43.75 52.92 43.838 ;
        RECT 35.946 43.796 52.874 43.884 ;
        RECT 35.9 43.842 52.828 43.93 ;
        RECT 35.854 43.888 52.782 43.976 ;
        RECT 35.808 43.934 52.736 44.022 ;
        RECT 35.762 43.98 52.69 44.068 ;
        RECT 35.716 44.026 52.644 44.114 ;
        RECT 35.67 44.072 52.598 44.16 ;
        RECT 35.624 44.118 52.552 44.206 ;
        RECT 35.578 44.164 52.506 44.252 ;
        RECT 35.532 44.21 52.46 44.298 ;
        RECT 35.486 44.256 52.414 44.344 ;
        RECT 35.44 44.302 52.368 44.39 ;
        RECT 35.394 44.348 52.322 44.436 ;
        RECT 35.348 44.394 52.276 44.482 ;
        RECT 35.302 44.44 52.23 44.528 ;
        RECT 35.256 44.486 52.184 44.574 ;
        RECT 35.21 44.532 52.138 44.62 ;
        RECT 35.164 44.578 52.092 44.666 ;
        RECT 35.118 44.624 52.046 44.712 ;
        RECT 35.072 44.67 52 44.758 ;
        RECT 35.026 44.716 51.954 44.804 ;
        RECT 34.98 44.762 51.908 44.85 ;
        RECT 34.934 44.808 51.862 44.896 ;
        RECT 34.888 44.854 51.816 44.942 ;
        RECT 34.842 44.9 51.77 44.988 ;
        RECT 34.796 44.946 51.724 45.034 ;
        RECT 34.75 44.992 51.678 45.08 ;
        RECT 34.704 45.038 51.632 45.126 ;
        RECT 34.658 45.084 51.586 45.172 ;
        RECT 34.612 45.13 51.54 45.218 ;
        RECT 34.566 45.176 51.494 45.264 ;
        RECT 34.52 45.222 51.448 45.31 ;
        RECT 34.474 45.268 51.402 45.356 ;
        RECT 34.428 45.314 51.356 45.402 ;
        RECT 34.382 45.36 51.31 45.448 ;
        RECT 34.336 45.406 51.264 45.494 ;
        RECT 34.29 45.452 51.218 45.54 ;
        RECT 34.244 45.498 51.172 45.586 ;
        RECT 34.198 45.544 51.126 45.632 ;
        RECT 34.152 45.59 51.08 45.678 ;
        RECT 34.106 45.636 51.034 45.724 ;
        RECT 34.06 45.682 50.988 45.77 ;
        RECT 34.014 45.728 50.942 45.816 ;
        RECT 33.968 45.774 50.896 45.862 ;
        RECT 33.922 45.82 50.85 45.908 ;
        RECT 33.876 45.866 50.804 45.954 ;
        RECT 33.83 45.912 50.758 46 ;
        RECT 33.784 45.958 50.712 46.046 ;
        RECT 33.738 46.004 50.666 46.092 ;
        RECT 33.692 46.05 50.62 46.138 ;
        RECT 33.646 46.096 50.574 46.184 ;
        RECT 33.6 46.142 50.528 46.23 ;
        RECT 33.554 46.188 50.482 46.276 ;
        RECT 33.508 46.234 50.436 46.322 ;
        RECT 33.462 46.28 50.39 46.368 ;
        RECT 33.416 46.326 50.344 46.414 ;
        RECT 33.37 46.372 50.298 46.46 ;
        RECT 33.324 46.418 50.252 46.506 ;
        RECT 33.278 46.464 50.206 46.552 ;
        RECT 33.232 46.51 50.16 46.598 ;
        RECT 33.186 46.556 50.114 46.644 ;
        RECT 33.14 46.602 50.068 46.69 ;
        RECT 33.094 46.648 50.022 46.736 ;
        RECT 33.048 46.694 49.976 46.782 ;
        RECT 33.002 46.74 49.93 46.828 ;
        RECT 32.956 46.786 49.884 46.874 ;
        RECT 32.91 46.832 49.838 46.92 ;
        RECT 32.864 46.878 49.792 46.966 ;
        RECT 32.818 46.924 49.746 47.012 ;
        RECT 32.772 46.97 49.7 47.058 ;
        RECT 32.726 47.016 49.654 47.104 ;
        RECT 32.68 47.062 49.608 47.15 ;
        RECT 32.634 47.108 49.562 47.196 ;
        RECT 32.588 47.154 49.516 47.242 ;
        RECT 32.542 47.2 49.47 47.288 ;
        RECT 32.496 47.246 49.424 47.334 ;
        RECT 32.45 47.292 49.378 47.38 ;
        RECT 32.404 47.338 49.332 47.426 ;
        RECT 32.358 47.384 49.286 47.472 ;
        RECT 32.312 47.43 49.24 47.518 ;
        RECT 32.266 47.476 49.194 47.564 ;
        RECT 32.22 47.522 49.148 47.61 ;
        RECT 32.174 47.568 49.102 47.656 ;
        RECT 32.128 47.614 49.056 47.702 ;
        RECT 32.082 47.66 49.01 47.748 ;
        RECT 32.036 47.706 48.964 47.794 ;
        RECT 31.99 47.752 48.918 47.84 ;
        RECT 31.944 47.798 48.872 47.886 ;
        RECT 31.898 47.844 48.826 47.932 ;
        RECT 31.852 47.89 48.78 47.978 ;
        RECT 31.806 47.936 48.734 48.024 ;
        RECT 31.76 47.982 48.688 48.07 ;
        RECT 31.714 48.028 48.642 48.116 ;
        RECT 31.668 48.074 48.596 48.162 ;
        RECT 31.622 48.12 48.55 48.208 ;
        RECT 31.576 48.166 48.504 48.254 ;
        RECT 31.53 48.212 48.458 48.3 ;
        RECT 31.484 48.258 48.412 48.346 ;
        RECT 31.438 48.304 48.366 48.392 ;
        RECT 31.392 48.35 48.32 48.438 ;
        RECT 31.346 48.396 48.274 48.484 ;
        RECT 31.3 48.442 48.228 48.53 ;
        RECT 31.254 48.488 48.182 48.576 ;
        RECT 31.208 48.534 48.136 48.622 ;
        RECT 31.162 48.58 48.09 48.668 ;
        RECT 31.116 48.626 48.044 48.714 ;
        RECT 31.07 48.672 47.998 48.76 ;
        RECT 31.024 48.718 47.952 48.806 ;
        RECT 30.978 48.764 47.906 48.852 ;
        RECT 30.932 48.81 47.86 48.898 ;
        RECT 30.886 48.856 47.814 48.944 ;
        RECT 30.84 48.902 47.768 48.99 ;
        RECT 30.794 48.948 47.722 49.036 ;
        RECT 30.748 48.994 47.676 49.082 ;
        RECT 30.702 49.04 47.63 49.128 ;
        RECT 30.656 49.086 47.584 49.174 ;
        RECT 30.61 49.132 47.538 49.22 ;
        RECT 30.564 49.178 47.492 49.266 ;
        RECT 30.518 49.224 47.446 49.312 ;
        RECT 30.472 49.27 47.4 49.358 ;
        RECT 30.426 49.316 47.354 49.404 ;
        RECT 30.38 49.362 47.308 49.45 ;
        RECT 30.334 49.408 47.262 49.496 ;
        RECT 30.288 49.454 47.216 49.542 ;
        RECT 30.242 49.5 47.17 49.588 ;
        RECT 30.196 49.546 47.124 49.634 ;
        RECT 30.15 49.592 47.078 49.68 ;
        RECT 30.104 49.638 47.032 49.726 ;
        RECT 30.058 49.684 46.986 49.772 ;
        RECT 30.012 49.73 46.94 49.818 ;
        RECT 29.966 49.776 46.894 49.864 ;
        RECT 29.92 49.822 46.848 49.91 ;
        RECT 29.874 49.868 46.802 49.956 ;
        RECT 29.828 49.914 46.756 50.002 ;
        RECT 29.782 49.96 46.71 50.048 ;
        RECT 29.736 50.006 46.664 50.094 ;
        RECT 29.69 50.052 46.618 50.14 ;
        RECT 29.644 50.098 46.572 50.186 ;
        RECT 29.598 50.144 46.526 50.232 ;
        RECT 29.552 50.19 46.48 50.278 ;
        RECT 29.506 50.236 46.434 50.324 ;
        RECT 29.46 50.282 46.388 50.37 ;
        RECT 29.414 50.328 46.342 50.416 ;
        RECT 29.368 50.374 46.296 50.462 ;
        RECT 29.322 50.42 46.25 50.508 ;
        RECT 29.276 50.466 46.204 50.554 ;
        RECT 29.23 50.512 46.158 50.6 ;
        RECT 29.184 50.558 46.112 50.646 ;
        RECT 29.138 50.604 46.066 50.692 ;
        RECT 29.092 50.65 46.02 50.738 ;
        RECT 29 50.742 45.974 50.784 ;
        RECT 29.046 50.696 45.974 50.784 ;
        RECT 28.96 50.785 45.928 50.83 ;
        RECT 28.914 50.828 45.882 50.876 ;
        RECT 28.868 50.874 45.836 50.922 ;
        RECT 28.822 50.92 45.79 50.968 ;
        RECT 28.776 50.966 45.744 51.014 ;
        RECT 28.73 51.012 45.698 51.06 ;
        RECT 28.684 51.058 45.652 51.106 ;
        RECT 28.638 51.104 45.606 51.152 ;
        RECT 28.592 51.15 45.56 51.198 ;
        RECT 28.546 51.196 45.514 51.244 ;
        RECT 28.5 51.242 45.468 51.29 ;
        RECT 28.454 51.288 45.422 51.336 ;
        RECT 28.408 51.334 45.376 51.382 ;
        RECT 56.015 3.5 110 15.5 ;
        RECT 39.052 20.44 56.015 20.488 ;
        RECT 39.098 20.394 56.061 20.447 ;
        RECT 55.98 3.517 56.015 20.488 ;
        RECT 39.144 20.348 56.107 20.401 ;
        RECT 55.934 3.558 55.98 20.528 ;
        RECT 39.006 20.486 55.934 20.574 ;
        RECT 39.19 20.302 56.153 20.355 ;
        RECT 55.888 3.604 55.934 20.574 ;
        RECT 38.96 20.532 55.888 20.62 ;
        RECT 39.236 20.256 56.199 20.309 ;
        RECT 55.842 3.65 55.888 20.62 ;
        RECT 38.914 20.578 55.842 20.666 ;
        RECT 39.282 20.21 56.245 20.263 ;
        RECT 55.796 3.696 55.842 20.666 ;
        RECT 38.868 20.624 55.796 20.712 ;
        RECT 39.328 20.164 56.291 20.217 ;
        RECT 55.75 3.742 55.796 20.712 ;
        RECT 38.822 20.67 55.75 20.758 ;
        RECT 39.374 20.118 56.337 20.171 ;
        RECT 55.704 3.788 55.75 20.758 ;
        RECT 38.776 20.716 55.704 20.804 ;
        RECT 39.42 20.072 56.383 20.125 ;
        RECT 55.658 3.834 55.704 20.804 ;
        RECT 38.73 20.762 55.658 20.85 ;
        RECT 39.466 20.026 56.429 20.079 ;
        RECT 55.612 3.88 55.658 20.85 ;
        RECT 38.684 20.808 55.612 20.896 ;
        RECT 39.512 19.98 56.475 20.033 ;
        RECT 55.566 3.926 55.612 20.896 ;
        RECT 38.638 20.854 55.566 20.942 ;
        RECT 39.558 19.934 56.521 19.987 ;
        RECT 55.52 3.972 55.566 20.942 ;
        RECT 38.592 20.9 55.52 20.988 ;
        RECT 39.604 19.888 56.567 19.941 ;
        RECT 55.474 4.018 55.52 20.988 ;
        RECT 38.546 20.946 55.474 21.034 ;
        RECT 39.65 19.842 56.613 19.895 ;
        RECT 55.428 4.064 55.474 21.034 ;
        RECT 38.5 20.992 55.428 21.08 ;
        RECT 39.696 19.796 56.659 19.849 ;
        RECT 55.382 4.11 55.428 21.08 ;
        RECT 38.454 21.038 55.382 21.126 ;
        RECT 39.742 19.75 56.705 19.803 ;
        RECT 55.336 4.156 55.382 21.126 ;
        RECT 38.408 21.084 55.336 21.172 ;
        RECT 39.788 19.704 56.751 19.757 ;
        RECT 55.29 4.202 55.336 21.172 ;
        RECT 38.362 21.13 55.29 21.218 ;
        RECT 39.834 19.658 56.797 19.711 ;
        RECT 55.244 4.248 55.29 21.218 ;
        RECT 38.316 21.176 55.244 21.264 ;
        RECT 39.88 19.612 56.843 19.665 ;
        RECT 55.198 4.294 55.244 21.264 ;
        RECT 38.27 21.222 55.198 21.31 ;
        RECT 39.926 19.566 56.889 19.619 ;
        RECT 55.152 4.34 55.198 21.31 ;
        RECT 38.224 21.268 55.152 21.356 ;
        RECT 39.972 19.52 56.935 19.573 ;
        RECT 55.106 4.386 55.152 21.356 ;
        RECT 38.178 21.314 55.106 21.402 ;
        RECT 40.018 19.474 56.981 19.527 ;
        RECT 55.06 4.432 55.106 21.402 ;
        RECT 38.132 21.36 55.06 21.448 ;
        RECT 40.064 19.428 57.027 19.481 ;
        RECT 55.014 4.478 55.06 21.448 ;
        RECT 38.086 21.406 55.014 21.494 ;
        RECT 40.11 19.382 57.073 19.435 ;
        RECT 54.968 4.524 55.014 21.494 ;
        RECT 38.04 21.452 54.968 21.54 ;
        RECT 40.156 19.336 57.119 19.389 ;
        RECT 54.922 4.57 54.968 21.54 ;
        RECT 37.994 21.498 54.922 21.586 ;
        RECT 40.202 19.29 57.165 19.343 ;
        RECT 54.876 4.616 54.922 21.586 ;
        RECT 37.948 21.544 54.876 21.632 ;
        RECT 40.248 19.244 57.211 19.297 ;
        RECT 54.83 4.662 54.876 21.632 ;
        RECT 37.902 21.59 54.83 21.678 ;
        RECT 40.294 19.198 57.257 19.251 ;
        RECT 54.784 4.708 54.83 21.678 ;
        RECT 37.856 21.636 54.784 21.724 ;
        RECT 40.34 19.152 57.303 19.205 ;
        RECT 54.738 4.754 54.784 21.724 ;
        RECT 37.81 21.682 54.738 21.77 ;
        RECT 40.386 19.106 57.349 19.159 ;
        RECT 54.692 4.8 54.738 21.77 ;
        RECT 37.764 21.728 54.692 21.816 ;
        RECT 40.432 19.06 57.395 19.113 ;
        RECT 54.646 4.846 54.692 21.816 ;
        RECT 37.718 21.774 54.646 21.862 ;
        RECT 40.478 19.014 57.441 19.067 ;
        RECT 54.6 4.892 54.646 21.862 ;
        RECT 37.672 21.82 54.6 21.908 ;
        RECT 40.524 18.968 57.487 19.021 ;
        RECT 54.554 4.938 54.6 21.908 ;
        RECT 37.626 21.866 54.554 21.954 ;
        RECT 40.57 18.922 57.533 18.975 ;
        RECT 54.508 4.984 54.554 21.954 ;
        RECT 37.58 21.912 54.508 22 ;
        RECT 40.616 18.876 57.579 18.929 ;
        RECT 54.462 5.03 54.508 22 ;
        RECT 37.534 21.958 54.462 22.046 ;
        RECT 40.662 18.83 57.625 18.883 ;
        RECT 54.416 5.076 54.462 22.046 ;
        RECT 37.488 22.004 54.416 22.092 ;
        RECT 40.708 18.784 57.671 18.837 ;
        RECT 54.37 5.122 54.416 22.092 ;
        RECT 37.442 22.05 54.37 22.138 ;
        RECT 40.754 18.738 57.717 18.791 ;
        RECT 54.324 5.168 54.37 22.138 ;
        RECT 37.396 22.096 54.324 22.184 ;
        RECT 40.8 18.692 57.763 18.745 ;
        RECT 54.278 5.214 54.324 22.184 ;
        RECT 37.35 22.142 54.278 22.23 ;
        RECT 40.846 18.646 57.809 18.699 ;
        RECT 54.232 5.26 54.278 22.23 ;
        RECT 37.304 22.188 54.232 22.276 ;
        RECT 40.892 18.6 57.855 18.653 ;
        RECT 54.186 5.306 54.232 22.276 ;
        RECT 37.258 22.234 54.186 22.322 ;
        RECT 40.938 18.554 57.901 18.607 ;
        RECT 54.14 5.352 54.186 22.322 ;
        RECT 37.212 22.28 54.14 22.368 ;
        RECT 40.984 18.508 57.947 18.561 ;
        RECT 54.094 5.398 54.14 22.368 ;
        RECT 37.166 22.326 54.094 22.414 ;
        RECT 41.03 18.462 57.993 18.515 ;
        RECT 54.048 5.444 54.094 22.414 ;
        RECT 37.12 22.372 54.048 22.46 ;
        RECT 41.076 18.416 58.039 18.469 ;
        RECT 54.002 5.49 54.048 22.46 ;
        RECT 37.074 22.418 54.002 22.506 ;
        RECT 41.122 18.37 58.085 18.423 ;
        RECT 53.956 5.536 54.002 22.506 ;
        RECT 37.028 22.464 53.956 22.552 ;
        RECT 41.168 18.324 58.131 18.377 ;
        RECT 53.91 5.582 53.956 22.552 ;
        RECT 36.982 22.51 53.91 22.598 ;
        RECT 41.214 18.278 58.177 18.331 ;
        RECT 53.864 5.628 53.91 22.598 ;
        RECT 36.936 22.556 53.864 22.644 ;
        RECT 41.26 18.232 58.223 18.285 ;
        RECT 53.818 5.674 53.864 22.644 ;
        RECT 36.89 22.602 53.818 22.69 ;
        RECT 41.306 18.186 58.269 18.239 ;
        RECT 53.772 5.72 53.818 22.69 ;
        RECT 36.844 22.648 53.772 22.736 ;
        RECT 41.352 18.14 58.315 18.193 ;
        RECT 53.726 5.766 53.772 22.736 ;
        RECT 36.798 22.694 53.726 22.782 ;
        RECT 41.398 18.094 58.361 18.147 ;
        RECT 53.68 5.812 53.726 22.782 ;
        RECT 36.752 22.74 53.68 22.828 ;
        RECT 41.444 18.048 58.407 18.101 ;
        RECT 53.634 5.858 53.68 22.828 ;
        RECT 36.706 22.786 53.634 22.874 ;
        RECT 41.49 18.002 58.453 18.055 ;
        RECT 53.588 5.904 53.634 22.874 ;
        RECT 36.66 22.832 53.588 22.92 ;
        RECT 41.536 17.956 58.499 18.009 ;
        RECT 53.542 5.95 53.588 22.92 ;
        RECT 36.614 22.878 53.542 22.966 ;
        RECT 41.582 17.91 58.545 17.963 ;
        RECT 53.496 5.996 53.542 22.966 ;
        RECT 36.568 22.924 53.496 23.012 ;
        RECT 41.628 17.864 58.591 17.917 ;
        RECT 53.45 6.042 53.496 23.012 ;
        RECT 36.522 22.97 53.45 23.058 ;
        RECT 41.674 17.818 58.637 17.871 ;
        RECT 53.404 6.088 53.45 23.058 ;
        RECT 36.476 23.016 53.404 23.104 ;
        RECT 41.72 17.772 58.683 17.825 ;
        RECT 53.358 6.134 53.404 23.104 ;
        RECT 36.43 23.062 53.358 23.15 ;
        RECT 41.766 17.726 58.729 17.779 ;
        RECT 53.312 6.18 53.358 23.15 ;
        RECT 36.384 23.108 53.312 23.196 ;
        RECT 41.812 17.68 58.775 17.733 ;
        RECT 53.266 6.226 53.312 23.196 ;
        RECT 36.338 23.154 53.266 23.242 ;
        RECT 41.858 17.634 58.821 17.687 ;
        RECT 53.22 6.272 53.266 23.242 ;
        RECT 36.292 23.2 53.22 23.288 ;
        RECT 41.904 17.588 58.867 17.641 ;
        RECT 53.174 6.318 53.22 23.288 ;
        RECT 36.246 23.246 53.174 23.334 ;
        RECT 41.95 17.542 58.913 17.595 ;
        RECT 53.128 6.364 53.174 23.334 ;
        RECT 36.2 23.292 53.128 23.38 ;
        RECT 41.996 17.496 58.959 17.549 ;
        RECT 53.082 6.41 53.128 23.38 ;
        RECT 36.154 23.338 53.082 23.426 ;
        RECT 42.042 17.45 59.005 17.503 ;
        RECT 53.036 6.456 53.082 23.426 ;
        RECT 36.108 23.384 53.036 23.472 ;
        RECT 42.088 17.404 59.051 17.457 ;
        RECT 52.99 6.502 53.036 23.472 ;
        RECT 36.062 23.43 52.99 23.518 ;
        RECT 42.134 17.358 59.097 17.411 ;
        RECT 52.944 6.548 52.99 23.518 ;
        RECT 36.016 23.476 52.944 23.564 ;
        RECT 42.18 17.312 59.143 17.365 ;
        RECT 52.898 6.594 52.944 23.564 ;
        RECT 35.97 23.522 52.898 23.61 ;
        RECT 42.226 17.266 59.189 17.319 ;
        RECT 52.852 6.64 52.898 23.61 ;
        RECT 35.924 23.568 52.852 23.656 ;
        RECT 42.272 17.22 59.235 17.273 ;
        RECT 52.806 6.686 52.852 23.656 ;
        RECT 35.878 23.614 52.806 23.702 ;
        RECT 42.318 17.174 59.281 17.227 ;
        RECT 52.76 6.732 52.806 23.702 ;
        RECT 35.832 23.66 52.76 23.748 ;
        RECT 42.364 17.128 59.327 17.181 ;
        RECT 52.714 6.778 52.76 23.748 ;
        RECT 35.786 23.706 52.714 23.794 ;
        RECT 42.41 17.082 59.373 17.135 ;
        RECT 52.668 6.824 52.714 23.794 ;
        RECT 35.74 23.752 52.668 23.84 ;
        RECT 42.456 17.036 59.419 17.089 ;
        RECT 52.622 6.87 52.668 23.84 ;
        RECT 35.694 23.798 52.622 23.886 ;
        RECT 42.502 16.99 59.465 17.043 ;
        RECT 52.576 6.916 52.622 23.886 ;
        RECT 35.648 23.844 52.576 23.932 ;
        RECT 42.548 16.944 59.511 16.997 ;
        RECT 52.53 6.962 52.576 23.932 ;
        RECT 35.602 23.89 52.53 23.978 ;
        RECT 42.594 16.898 59.557 16.951 ;
        RECT 52.484 7.008 52.53 23.978 ;
        RECT 35.556 23.936 52.484 24.024 ;
        RECT 42.64 16.852 59.603 16.905 ;
        RECT 52.438 7.054 52.484 24.024 ;
        RECT 35.51 23.982 52.438 24.07 ;
        RECT 42.686 16.806 59.649 16.859 ;
        RECT 52.392 7.1 52.438 24.07 ;
        RECT 35.464 24.028 52.392 24.116 ;
        RECT 42.732 16.76 59.695 16.813 ;
        RECT 52.346 7.146 52.392 24.116 ;
        RECT 35.418 24.074 52.346 24.162 ;
        RECT 42.778 16.714 59.741 16.767 ;
        RECT 52.3 7.192 52.346 24.162 ;
        RECT 35.372 24.12 52.3 24.208 ;
        RECT 42.824 16.668 59.787 16.721 ;
        RECT 52.254 7.238 52.3 24.208 ;
        RECT 35.326 24.166 52.254 24.254 ;
        RECT 42.87 16.622 59.833 16.675 ;
        RECT 52.208 7.284 52.254 24.254 ;
        RECT 35.28 24.212 52.208 24.3 ;
        RECT 42.916 16.576 59.879 16.629 ;
        RECT 52.162 7.33 52.208 24.3 ;
        RECT 35.234 24.258 52.162 24.346 ;
        RECT 42.962 16.53 59.925 16.583 ;
        RECT 52.116 7.376 52.162 24.346 ;
        RECT 35.188 24.304 52.116 24.392 ;
        RECT 43.008 16.484 59.971 16.537 ;
        RECT 52.07 7.422 52.116 24.392 ;
        RECT 35.142 24.35 52.07 24.438 ;
        RECT 43.054 16.438 60.017 16.491 ;
        RECT 52.024 7.468 52.07 24.438 ;
        RECT 35.096 24.396 52.024 24.484 ;
        RECT 43.1 16.392 60.063 16.445 ;
        RECT 51.978 7.514 52.024 24.484 ;
        RECT 35.05 24.442 51.978 24.53 ;
        RECT 43.146 16.346 60.109 16.399 ;
        RECT 51.932 7.56 51.978 24.53 ;
        RECT 35.004 24.488 51.932 24.576 ;
        RECT 43.192 16.3 60.155 16.353 ;
        RECT 51.886 7.606 51.932 24.576 ;
        RECT 34.958 24.534 51.886 24.622 ;
        RECT 43.238 16.254 60.201 16.307 ;
        RECT 51.84 7.652 51.886 24.622 ;
        RECT 34.912 24.58 51.84 24.668 ;
        RECT 43.284 16.208 60.247 16.261 ;
        RECT 51.794 7.698 51.84 24.668 ;
        RECT 34.866 24.626 51.794 24.714 ;
        RECT 43.33 16.162 60.293 16.215 ;
        RECT 51.748 7.744 51.794 24.714 ;
        RECT 34.82 24.672 51.748 24.76 ;
        RECT 43.376 16.116 60.339 16.169 ;
        RECT 51.702 7.79 51.748 24.76 ;
        RECT 34.774 24.718 51.702 24.806 ;
        RECT 43.422 16.07 60.385 16.123 ;
        RECT 51.656 7.836 51.702 24.806 ;
        RECT 34.728 24.764 51.656 24.852 ;
        RECT 43.468 16.024 60.431 16.077 ;
        RECT 51.61 7.882 51.656 24.852 ;
        RECT 34.682 24.81 51.61 24.898 ;
        RECT 43.514 15.978 60.477 16.031 ;
        RECT 51.564 7.928 51.61 24.898 ;
        RECT 34.636 24.856 51.564 24.944 ;
        RECT 43.56 15.932 60.523 15.985 ;
        RECT 51.518 7.974 51.564 24.944 ;
        RECT 34.59 24.902 51.518 24.99 ;
        RECT 43.606 15.886 60.569 15.939 ;
        RECT 51.472 8.02 51.518 24.99 ;
        RECT 34.544 24.948 51.472 25.036 ;
        RECT 43.652 15.84 60.615 15.893 ;
        RECT 51.426 8.066 51.472 25.036 ;
        RECT 34.498 24.994 51.426 25.082 ;
        RECT 43.698 15.794 60.661 15.847 ;
        RECT 51.38 8.112 51.426 25.082 ;
        RECT 34.452 25.04 51.38 25.128 ;
        RECT 43.744 15.748 60.707 15.801 ;
        RECT 51.334 8.158 51.38 25.128 ;
        RECT 34.406 25.086 51.334 25.174 ;
        RECT 43.79 15.702 60.753 15.755 ;
        RECT 51.288 8.204 51.334 25.174 ;
        RECT 34.36 25.132 51.288 25.22 ;
        RECT 43.836 15.656 60.799 15.709 ;
        RECT 51.242 8.25 51.288 25.22 ;
        RECT 34.314 25.178 51.242 25.266 ;
        RECT 43.882 15.61 60.845 15.663 ;
        RECT 51.196 8.296 51.242 25.266 ;
        RECT 34.268 25.224 51.196 25.312 ;
        RECT 43.928 15.564 60.891 15.617 ;
        RECT 51.15 8.342 51.196 25.312 ;
        RECT 34.222 25.27 51.15 25.358 ;
        RECT 43.974 15.518 60.937 15.571 ;
        RECT 51.104 8.388 51.15 25.358 ;
        RECT 34.176 25.316 51.104 25.404 ;
        RECT 44.02 15.472 60.983 15.524 ;
        RECT 51.058 8.434 51.104 25.404 ;
        RECT 34.13 25.362 51.058 25.45 ;
        RECT 44.066 15.426 110 15.5 ;
        RECT 51.012 8.48 51.058 25.45 ;
        RECT 34.084 25.408 51.012 25.496 ;
        RECT 44.112 15.38 110 15.5 ;
        RECT 50.966 8.526 51.012 25.496 ;
        RECT 34.038 25.454 50.966 25.542 ;
        RECT 44.158 15.334 110 15.5 ;
        RECT 50.92 8.572 50.966 25.542 ;
        RECT 33.992 25.5 50.92 25.588 ;
        RECT 44.204 15.288 110 15.5 ;
        RECT 50.874 8.618 50.92 25.588 ;
        RECT 33.946 25.546 50.874 25.634 ;
        RECT 44.25 15.242 110 15.5 ;
        RECT 50.828 8.664 50.874 25.634 ;
        RECT 33.9 25.592 50.828 25.68 ;
        RECT 44.296 15.196 110 15.5 ;
        RECT 50.782 8.71 50.828 25.68 ;
        RECT 33.854 25.638 50.782 25.726 ;
        RECT 44.342 15.15 110 15.5 ;
        RECT 50.736 8.756 50.782 25.726 ;
        RECT 33.808 25.684 50.736 25.772 ;
        RECT 44.388 15.104 110 15.5 ;
        RECT 50.69 8.802 50.736 25.772 ;
        RECT 33.762 25.73 50.69 25.818 ;
        RECT 44.434 15.058 110 15.5 ;
        RECT 50.644 8.848 50.69 25.818 ;
        RECT 33.716 25.776 50.644 25.864 ;
        RECT 44.48 15.012 110 15.5 ;
        RECT 50.598 8.894 50.644 25.864 ;
        RECT 33.67 25.822 50.598 25.91 ;
        RECT 44.526 14.966 110 15.5 ;
        RECT 50.552 8.94 50.598 25.91 ;
        RECT 33.624 25.868 50.552 25.956 ;
        RECT 44.572 14.92 110 15.5 ;
        RECT 50.506 8.986 50.552 25.956 ;
        RECT 33.578 25.914 50.506 26.002 ;
        RECT 44.618 14.874 110 15.5 ;
        RECT 50.46 9.032 50.506 26.002 ;
        RECT 33.532 25.96 50.46 26.048 ;
        RECT 44.664 14.828 110 15.5 ;
        RECT 50.414 9.078 50.46 26.048 ;
        RECT 33.486 26.006 50.414 26.094 ;
        RECT 44.71 14.782 110 15.5 ;
        RECT 50.368 9.124 50.414 26.094 ;
        RECT 33.44 26.052 50.368 26.14 ;
        RECT 44.756 14.736 110 15.5 ;
        RECT 50.322 9.17 50.368 26.14 ;
        RECT 33.394 26.098 50.322 26.186 ;
        RECT 44.802 14.69 110 15.5 ;
        RECT 50.276 9.216 50.322 26.186 ;
        RECT 33.348 26.144 50.276 26.232 ;
        RECT 44.848 14.644 110 15.5 ;
        RECT 50.23 9.262 50.276 26.232 ;
        RECT 33.302 26.19 50.23 26.278 ;
        RECT 44.894 14.598 110 15.5 ;
        RECT 50.184 9.308 50.23 26.278 ;
        RECT 33.256 26.236 50.184 26.324 ;
        RECT 44.94 14.552 110 15.5 ;
        RECT 50.138 9.354 50.184 26.324 ;
        RECT 33.21 26.282 50.138 26.37 ;
        RECT 44.986 14.506 110 15.5 ;
        RECT 50.092 9.4 50.138 26.37 ;
        RECT 33.164 26.328 50.092 26.416 ;
        RECT 45.032 14.46 110 15.5 ;
        RECT 50.046 9.446 50.092 26.416 ;
        RECT 33.118 26.374 50.046 26.462 ;
        RECT 45.078 14.414 110 15.5 ;
        RECT 50 9.492 50.046 26.462 ;
        RECT 33.072 26.42 50 26.508 ;
        RECT 45.124 14.368 110 15.5 ;
        RECT 49.954 9.538 50 26.508 ;
        RECT 33.026 26.466 49.954 26.554 ;
        RECT 45.17 14.322 110 15.5 ;
        RECT 49.908 9.584 49.954 26.554 ;
        RECT 32.98 26.512 49.908 26.6 ;
        RECT 45.216 14.276 110 15.5 ;
        RECT 49.862 9.63 49.908 26.6 ;
        RECT 32.934 26.558 49.862 26.646 ;
        RECT 45.262 14.23 110 15.5 ;
        RECT 49.816 9.676 49.862 26.646 ;
        RECT 32.888 26.604 49.816 26.692 ;
        RECT 45.308 14.184 110 15.5 ;
        RECT 49.77 9.722 49.816 26.692 ;
        RECT 32.842 26.65 49.77 26.738 ;
        RECT 45.354 14.138 110 15.5 ;
        RECT 49.724 9.768 49.77 26.738 ;
        RECT 32.796 26.696 49.724 26.784 ;
        RECT 45.4 14.092 110 15.5 ;
        RECT 49.678 9.814 49.724 26.784 ;
        RECT 32.75 26.742 49.678 26.83 ;
        RECT 45.446 14.046 110 15.5 ;
        RECT 49.632 9.86 49.678 26.83 ;
        RECT 32.704 26.788 49.632 26.876 ;
        RECT 45.492 14 110 15.5 ;
        RECT 49.586 9.906 49.632 26.876 ;
        RECT 32.658 26.834 49.586 26.922 ;
        RECT 45.538 13.954 110 15.5 ;
        RECT 49.54 9.952 49.586 26.922 ;
        RECT 32.612 26.88 49.54 26.968 ;
        RECT 45.584 13.908 110 15.5 ;
        RECT 49.494 9.998 49.54 26.968 ;
        RECT 32.566 26.926 49.494 27.014 ;
        RECT 45.63 13.862 110 15.5 ;
        RECT 49.448 10.044 49.494 27.014 ;
        RECT 32.52 26.972 49.448 27.06 ;
        RECT 45.676 13.816 110 15.5 ;
        RECT 49.402 10.09 49.448 27.06 ;
        RECT 32.474 27.018 49.402 27.106 ;
        RECT 45.722 13.77 110 15.5 ;
        RECT 49.356 10.136 49.402 27.106 ;
        RECT 32.428 27.064 49.356 27.152 ;
        RECT 45.768 13.724 110 15.5 ;
        RECT 49.31 10.182 49.356 27.152 ;
        RECT 32.382 27.11 49.31 27.198 ;
        RECT 45.814 13.678 110 15.5 ;
        RECT 49.264 10.228 49.31 27.198 ;
        RECT 32.336 27.156 49.264 27.244 ;
        RECT 45.86 13.632 110 15.5 ;
        RECT 49.218 10.274 49.264 27.244 ;
        RECT 32.29 27.202 49.218 27.29 ;
        RECT 45.906 13.586 110 15.5 ;
        RECT 49.172 10.32 49.218 27.29 ;
        RECT 32.244 27.248 49.172 27.336 ;
        RECT 45.952 13.54 110 15.5 ;
        RECT 49.126 10.366 49.172 27.336 ;
        RECT 32.198 27.294 49.126 27.382 ;
        RECT 45.998 13.494 110 15.5 ;
        RECT 49.08 10.412 49.126 27.382 ;
        RECT 32.152 27.34 49.08 27.428 ;
        RECT 46.044 13.448 110 15.5 ;
        RECT 49.034 10.458 49.08 27.428 ;
        RECT 32.106 27.386 49.034 27.474 ;
        RECT 46.09 13.402 110 15.5 ;
        RECT 48.988 10.504 49.034 27.474 ;
        RECT 32.06 27.432 48.988 27.52 ;
        RECT 46.136 13.356 110 15.5 ;
        RECT 48.942 10.55 48.988 27.52 ;
        RECT 32.014 27.478 48.942 27.566 ;
        RECT 46.182 13.31 110 15.5 ;
        RECT 48.896 10.596 48.942 27.566 ;
        RECT 31.968 27.524 48.896 27.612 ;
        RECT 46.228 13.264 110 15.5 ;
        RECT 48.85 10.642 48.896 27.612 ;
        RECT 31.922 27.57 48.85 27.658 ;
        RECT 46.274 13.218 110 15.5 ;
        RECT 48.804 10.688 48.85 27.658 ;
        RECT 31.876 27.616 48.804 27.704 ;
        RECT 46.32 13.172 110 15.5 ;
        RECT 48.758 10.734 48.804 27.704 ;
        RECT 31.83 27.662 48.758 27.75 ;
        RECT 46.366 13.126 110 15.5 ;
        RECT 48.712 10.78 48.758 27.75 ;
        RECT 31.784 27.708 48.712 27.796 ;
        RECT 46.412 13.08 110 15.5 ;
        RECT 48.666 10.826 48.712 27.796 ;
        RECT 31.738 27.754 48.666 27.842 ;
        RECT 46.458 13.034 110 15.5 ;
        RECT 48.62 10.872 48.666 27.842 ;
        RECT 31.692 27.8 48.62 27.888 ;
        RECT 46.504 12.988 110 15.5 ;
        RECT 48.574 10.918 48.62 27.888 ;
        RECT 31.646 27.846 48.574 27.934 ;
        RECT 46.55 12.942 110 15.5 ;
        RECT 48.528 10.964 48.574 27.934 ;
        RECT 31.6 27.892 48.528 27.98 ;
        RECT 46.596 12.896 110 15.5 ;
        RECT 48.482 11.01 48.528 27.98 ;
        RECT 31.554 27.938 48.482 28.026 ;
        RECT 46.642 12.85 110 15.5 ;
        RECT 48.436 11.056 48.482 28.026 ;
        RECT 31.508 27.984 48.436 28.072 ;
        RECT 46.688 12.804 110 15.5 ;
        RECT 48.39 11.102 48.436 28.072 ;
        RECT 31.462 28.03 48.39 28.118 ;
        RECT 46.734 12.758 110 15.5 ;
        RECT 48.344 11.148 48.39 28.118 ;
        RECT 31.416 28.076 48.344 28.164 ;
        RECT 46.78 12.712 110 15.5 ;
        RECT 48.298 11.194 48.344 28.164 ;
        RECT 31.37 28.122 48.298 28.21 ;
        RECT 46.826 12.666 110 15.5 ;
        RECT 48.252 11.24 48.298 28.21 ;
        RECT 31.324 28.168 48.252 28.256 ;
        RECT 46.872 12.62 110 15.5 ;
        RECT 48.206 11.286 48.252 28.256 ;
        RECT 31.278 28.214 48.206 28.302 ;
        RECT 46.918 12.574 110 15.5 ;
        RECT 48.16 11.332 48.206 28.302 ;
        RECT 31.232 28.26 48.16 28.348 ;
        RECT 46.964 12.528 110 15.5 ;
        RECT 48.114 11.378 48.16 28.348 ;
        RECT 31.186 28.306 48.114 28.394 ;
        RECT 47.01 12.482 110 15.5 ;
        RECT 48.068 11.424 48.114 28.394 ;
        RECT 31.14 28.352 48.068 28.44 ;
        RECT 47.056 12.436 110 15.5 ;
        RECT 48.022 11.47 48.068 28.44 ;
        RECT 31.094 28.398 48.022 28.486 ;
        RECT 47.102 12.39 110 15.5 ;
        RECT 47.976 11.516 48.022 28.486 ;
        RECT 31.048 28.444 47.976 28.532 ;
        RECT 47.148 12.344 110 15.5 ;
        RECT 47.93 11.562 47.976 28.532 ;
        RECT 31.002 28.49 47.93 28.578 ;
        RECT 47.194 12.298 110 15.5 ;
        RECT 47.884 11.608 47.93 28.578 ;
        RECT 30.956 28.536 47.884 28.624 ;
        RECT 47.24 12.252 110 15.5 ;
        RECT 47.838 11.654 47.884 28.624 ;
        RECT 30.91 28.582 47.838 28.67 ;
        RECT 47.286 12.206 110 15.5 ;
        RECT 47.792 11.7 47.838 28.67 ;
        RECT 30.864 28.628 47.792 28.716 ;
        RECT 47.332 12.16 110 15.5 ;
        RECT 47.746 11.746 47.792 28.716 ;
        RECT 30.818 28.674 47.746 28.762 ;
        RECT 47.378 12.114 110 15.5 ;
        RECT 47.7 11.792 47.746 28.762 ;
        RECT 30.772 28.72 47.7 28.808 ;
        RECT 47.424 12.068 110 15.5 ;
        RECT 47.654 11.838 47.7 28.808 ;
        RECT 30.726 28.766 47.654 28.854 ;
        RECT 47.47 12.022 110 15.5 ;
        RECT 47.608 11.884 47.654 28.854 ;
        RECT 30.68 28.812 47.608 28.9 ;
        RECT 47.516 11.976 110 15.5 ;
        RECT 47.562 11.93 47.608 28.9 ;
        RECT 30.634 28.858 47.562 28.946 ;
        RECT 30.588 28.904 47.516 28.992 ;
        RECT 30.542 28.95 47.47 29.038 ;
        RECT 30.496 28.996 47.424 29.084 ;
        RECT 30.45 29.042 47.378 29.13 ;
        RECT 30.404 29.088 47.332 29.176 ;
        RECT 30.358 29.134 47.286 29.222 ;
        RECT 30.312 29.18 47.24 29.268 ;
        RECT 30.266 29.226 47.194 29.314 ;
        RECT 30.22 29.272 47.148 29.36 ;
        RECT 30.174 29.318 47.102 29.406 ;
        RECT 30.128 29.364 47.056 29.452 ;
        RECT 30.082 29.41 47.01 29.498 ;
        RECT 30.036 29.456 46.964 29.544 ;
        RECT 29.99 29.502 46.918 29.59 ;
        RECT 29.944 29.548 46.872 29.636 ;
        RECT 29.898 29.594 46.826 29.682 ;
        RECT 29.852 29.64 46.78 29.728 ;
        RECT 29.806 29.686 46.734 29.774 ;
        RECT 29.76 29.732 46.688 29.82 ;
        RECT 29.714 29.778 46.642 29.866 ;
        RECT 29.668 29.824 46.596 29.912 ;
        RECT 29.622 29.87 46.55 29.958 ;
        RECT 29.576 29.916 46.504 30.004 ;
        RECT 29.53 29.962 46.458 30.05 ;
        RECT 29.484 30.008 46.412 30.096 ;
        RECT 29.438 30.054 46.366 30.142 ;
        RECT 29.392 30.1 46.32 30.188 ;
        RECT 29.346 30.146 46.274 30.234 ;
        RECT 29.3 30.192 46.228 30.28 ;
        RECT 29.254 30.238 46.182 30.326 ;
        RECT 29.208 30.284 46.136 30.372 ;
        RECT 29.162 30.33 46.09 30.418 ;
        RECT 29.116 30.376 46.044 30.464 ;
        RECT 29.07 30.422 45.998 30.51 ;
        RECT 29.024 30.468 45.952 30.556 ;
        RECT 28.978 30.514 45.906 30.602 ;
        RECT 28.932 30.56 45.86 30.648 ;
        RECT 28.886 30.606 45.814 30.694 ;
        RECT 28.84 30.652 45.768 30.74 ;
        RECT 28.794 30.698 45.722 30.786 ;
        RECT 28.748 30.744 45.676 30.832 ;
        RECT 28.702 30.79 45.63 30.878 ;
        RECT 28.656 30.836 45.584 30.924 ;
        RECT 28.61 30.882 45.538 30.97 ;
        RECT 28.564 30.928 45.492 31.016 ;
        RECT 28.518 30.974 45.446 31.062 ;
        RECT 28.472 31.02 45.4 31.108 ;
        RECT 28.426 31.066 45.354 31.154 ;
        RECT 28.38 31.112 45.308 31.2 ;
        RECT 28.334 31.158 45.262 31.246 ;
        RECT 28.288 31.204 45.216 31.292 ;
        RECT 28.242 31.25 45.17 31.338 ;
        RECT 28.196 31.296 45.124 31.384 ;
        RECT 28.15 31.342 45.078 31.43 ;
        RECT 28.104 31.388 45.032 31.476 ;
        RECT 28.058 31.434 44.986 31.522 ;
        RECT 28.012 31.48 44.94 31.568 ;
        RECT 27.966 31.526 44.894 31.614 ;
        RECT 27.92 31.572 44.848 31.66 ;
        RECT 27.874 31.618 44.802 31.706 ;
        RECT 27.828 31.664 44.756 31.752 ;
        RECT 27.782 31.71 44.71 31.798 ;
        RECT 27.736 31.756 44.664 31.844 ;
        RECT 27.69 31.802 44.618 31.89 ;
        RECT 27.644 31.848 44.572 31.936 ;
        RECT 27.598 31.894 44.526 31.982 ;
        RECT 27.552 31.94 44.48 32.028 ;
        RECT 27.506 31.986 44.434 32.074 ;
        RECT 27.46 32.032 44.388 32.12 ;
        RECT 27.414 32.078 44.342 32.166 ;
        RECT 27.368 32.124 44.296 32.212 ;
        RECT 27.322 32.17 44.25 32.258 ;
        RECT 27.276 32.216 44.204 32.304 ;
        RECT 27.23 32.262 44.158 32.35 ;
        RECT 27.184 32.308 44.112 32.396 ;
        RECT 27.138 32.354 44.066 32.442 ;
        RECT 27.092 32.4 44.02 32.488 ;
        RECT 27.046 32.446 43.974 32.534 ;
        RECT 27 32.492 43.928 32.58 ;
        RECT 26.954 32.538 43.882 32.626 ;
        RECT 26.908 32.584 43.836 32.672 ;
        RECT 26.862 32.63 43.79 32.718 ;
        RECT 26.816 32.676 43.744 32.764 ;
        RECT 26.77 32.722 43.698 32.81 ;
        RECT 26.724 32.768 43.652 32.856 ;
        RECT 26.678 32.814 43.606 32.902 ;
        RECT 26.632 32.86 43.56 32.948 ;
        RECT 26.586 32.906 43.514 32.994 ;
        RECT 26.54 32.952 43.468 33.04 ;
        RECT 26.494 32.998 43.422 33.086 ;
        RECT 26.448 33.044 43.376 33.132 ;
        RECT 26.402 33.09 43.33 33.178 ;
        RECT 26.356 33.136 43.284 33.224 ;
        RECT 26.31 33.182 43.238 33.27 ;
        RECT 26.264 33.228 43.192 33.316 ;
        RECT 26.218 33.274 43.146 33.362 ;
        RECT 26.172 33.32 43.1 33.408 ;
        RECT 26.126 33.366 43.054 33.454 ;
        RECT 26.08 33.412 43.008 33.5 ;
        RECT 26.034 33.458 42.962 33.546 ;
        RECT 25.988 33.504 42.916 33.592 ;
        RECT 25.942 33.55 42.87 33.638 ;
        RECT 25.896 33.596 42.824 33.684 ;
        RECT 25.85 33.642 42.778 33.73 ;
        RECT 25.804 33.688 42.732 33.776 ;
        RECT 25.758 33.734 42.686 33.822 ;
        RECT 25.712 33.78 42.64 33.868 ;
        RECT 25.666 33.826 42.594 33.914 ;
        RECT 25.62 33.872 42.548 33.96 ;
        RECT 25.574 33.918 42.502 34.006 ;
        RECT 25.528 33.964 42.456 34.052 ;
        RECT 25.482 34.01 42.41 34.098 ;
        RECT 25.436 34.056 42.364 34.144 ;
        RECT 25.39 34.102 42.318 34.19 ;
        RECT 25.344 34.148 42.272 34.236 ;
        RECT 25.298 34.194 42.226 34.282 ;
        RECT 25.252 34.24 42.18 34.328 ;
        RECT 25.206 34.286 42.134 34.374 ;
        RECT 25.16 34.332 42.088 34.42 ;
        RECT 25.114 34.378 42.042 34.466 ;
        RECT 25.068 34.424 41.996 34.512 ;
        RECT 25.022 34.47 41.95 34.558 ;
        RECT 24.976 34.516 41.904 34.604 ;
        RECT 24.93 34.562 41.858 34.65 ;
        RECT 24.884 34.608 41.812 34.696 ;
        RECT 24.838 34.654 41.766 34.742 ;
        RECT 24.792 34.7 41.72 34.788 ;
        RECT 24.746 34.746 41.674 34.834 ;
        RECT 24.7 34.792 41.628 34.88 ;
        RECT 24.654 34.838 41.582 34.926 ;
        RECT 24.608 34.884 41.536 34.972 ;
        RECT 24.562 34.93 41.49 35.018 ;
        RECT 24.516 34.976 41.444 35.064 ;
        RECT 24.47 35.022 41.398 35.11 ;
        RECT 24.424 35.068 41.352 35.156 ;
        RECT 24.378 35.114 41.306 35.202 ;
        RECT 24.332 35.16 41.26 35.248 ;
        RECT 24.286 35.206 41.214 35.294 ;
        RECT 24.24 35.252 41.168 35.34 ;
        RECT 24.194 35.298 41.122 35.386 ;
        RECT 24.148 35.344 41.076 35.432 ;
        RECT 24.102 35.39 41.03 35.478 ;
        RECT 24.056 35.436 40.984 35.524 ;
        RECT 24.01 35.482 40.938 35.57 ;
        RECT 23.964 35.528 40.892 35.616 ;
        RECT 23.918 35.574 40.846 35.662 ;
        RECT 23.872 35.62 40.8 35.708 ;
        RECT 23.826 35.666 40.754 35.754 ;
        RECT 23.78 35.712 40.708 35.8 ;
        RECT 23.734 35.758 40.662 35.846 ;
        RECT 23.688 35.804 40.616 35.892 ;
        RECT 23.642 35.85 40.57 35.938 ;
        RECT 23.596 35.896 40.524 35.984 ;
        RECT 23.55 35.942 40.478 36.03 ;
        RECT 23.504 35.988 40.432 36.076 ;
        RECT 23.458 36.034 40.386 36.122 ;
        RECT 23.412 36.08 40.34 36.168 ;
        RECT 23.366 36.126 40.294 36.214 ;
        RECT 23.32 36.172 40.248 36.26 ;
        RECT 23.274 36.218 40.202 36.306 ;
        RECT 23.228 36.264 40.156 36.352 ;
        RECT 23.182 36.31 40.11 36.398 ;
        RECT 23.136 36.356 40.064 36.444 ;
        RECT 23.09 36.402 40.018 36.49 ;
        RECT 23.044 36.448 39.972 36.536 ;
        RECT 22.998 36.494 39.926 36.582 ;
        RECT 22.952 36.54 39.88 36.628 ;
        RECT 22.906 36.586 39.834 36.674 ;
        RECT 22.86 36.632 39.788 36.72 ;
        RECT 22.814 36.678 39.742 36.766 ;
        RECT 22.768 36.724 39.696 36.812 ;
        RECT 22.722 36.77 39.65 36.858 ;
        RECT 22.676 36.816 39.604 36.904 ;
        RECT 22.63 36.862 39.558 36.95 ;
        RECT 22.584 36.908 39.512 36.996 ;
        RECT 22.538 36.954 39.466 37.042 ;
        RECT 22.492 37 39.42 37.088 ;
        RECT 22.446 37.046 39.374 37.134 ;
        RECT 22.4 37.092 39.328 37.18 ;
        RECT 22.354 37.138 39.282 37.226 ;
        RECT 22.308 37.184 39.236 37.272 ;
        RECT 22.262 37.23 39.19 37.318 ;
        RECT 22.216 37.276 39.144 37.364 ;
        RECT 22.17 37.322 39.098 37.41 ;
        RECT 22.124 37.368 39.052 37.456 ;
        RECT 22.078 37.414 39.006 37.502 ;
        RECT 22.032 37.46 38.96 37.548 ;
        RECT 21.986 37.506 38.914 37.594 ;
        RECT 21.94 37.552 38.868 37.64 ;
        RECT 21.894 37.598 38.822 37.686 ;
        RECT 21.848 37.644 38.776 37.732 ;
        RECT 21.802 37.69 38.73 37.778 ;
        RECT 21.756 37.736 38.684 37.824 ;
        RECT 21.71 37.782 38.638 37.87 ;
        RECT 21.664 37.828 38.592 37.916 ;
        RECT 21.618 37.874 38.546 37.962 ;
        RECT 21.572 37.92 38.5 38.008 ;
        RECT 21.526 37.966 38.454 38.054 ;
        RECT 21.48 38.012 38.408 38.1 ;
        RECT 21.434 38.058 38.362 38.146 ;
        RECT 21.388 38.104 38.316 38.192 ;
        RECT 21.342 38.15 38.27 38.238 ;
        RECT 21.296 38.196 38.224 38.284 ;
        RECT 21.25 38.242 38.178 38.33 ;
        RECT 21.204 38.288 38.132 38.376 ;
        RECT 21.158 38.334 38.086 38.422 ;
        RECT 21.112 38.38 38.04 38.468 ;
        RECT 21.066 38.426 37.994 38.514 ;
        RECT 21.02 38.472 37.948 38.56 ;
        RECT 20.974 38.518 37.902 38.606 ;
        RECT 20.928 38.564 37.856 38.652 ;
        RECT 20.882 38.61 37.81 38.698 ;
        RECT 20.836 38.656 37.764 38.744 ;
        RECT 20.79 38.702 37.718 38.79 ;
        RECT 20.744 38.748 37.672 38.836 ;
        RECT 20.698 38.794 37.626 38.882 ;
        RECT 20.652 38.84 37.58 38.928 ;
        RECT 20.606 38.886 37.534 38.974 ;
        RECT 20.56 38.932 37.488 39.02 ;
        RECT 20.514 38.978 37.442 39.066 ;
        RECT 20.468 39.024 37.396 39.112 ;
        RECT 20.422 39.07 37.35 39.158 ;
        RECT 20.376 39.116 37.304 39.204 ;
        RECT 20.33 39.162 37.258 39.25 ;
        RECT 20.284 39.208 37.212 39.296 ;
        RECT 20.238 39.254 37.166 39.342 ;
        RECT 20.192 39.3 37.12 39.388 ;
        RECT 20.146 39.346 37.074 39.434 ;
        RECT 20.1 39.392 37.028 39.48 ;
        RECT 20.054 39.438 36.982 39.526 ;
        RECT 20.008 39.484 36.936 39.572 ;
        RECT 19.962 39.53 36.89 39.618 ;
        RECT 19.916 39.576 36.844 39.664 ;
        RECT 19.87 39.622 36.798 39.71 ;
        RECT 19.824 39.668 36.752 39.756 ;
        RECT 19.778 39.714 36.706 39.802 ;
        RECT 19.732 39.76 36.66 39.848 ;
        RECT 19.686 39.806 36.614 39.894 ;
        RECT 19.64 39.852 36.568 39.94 ;
        RECT 19.594 39.898 36.522 39.986 ;
        RECT 19.548 39.944 36.476 40.032 ;
        RECT 19.502 39.99 36.43 40.078 ;
        RECT 19.456 40.036 36.384 40.124 ;
        RECT 19.41 40.082 36.338 40.17 ;
        RECT 19.364 40.128 36.292 40.216 ;
        RECT 19.318 40.174 36.246 40.262 ;
        RECT 19.272 40.22 36.2 40.308 ;
        RECT 19.226 40.266 36.154 40.354 ;
        RECT 19.18 40.312 36.108 40.4 ;
        RECT 19.134 40.358 36.062 40.446 ;
        RECT 19.088 40.404 36.016 40.492 ;
        RECT 19.042 40.45 35.97 40.538 ;
        RECT 18.996 40.496 35.924 40.584 ;
        RECT 18.95 40.542 35.878 40.63 ;
        RECT 18.904 40.588 35.832 40.676 ;
        RECT 18.858 40.634 35.786 40.722 ;
        RECT 18.812 40.68 35.74 40.768 ;
        RECT 18.766 40.726 35.694 40.814 ;
        RECT 18.72 40.772 35.648 40.86 ;
        RECT 18.674 40.818 35.602 40.906 ;
        RECT 18.628 40.864 35.556 40.952 ;
        RECT 18.582 40.91 35.51 40.998 ;
        RECT 18.536 40.956 35.464 41.044 ;
        RECT 18.49 41.002 35.418 41.09 ;
        RECT 18.444 41.048 35.372 41.136 ;
        RECT 18.398 41.094 35.326 41.182 ;
        RECT 18.352 41.14 35.28 41.228 ;
        RECT 18.306 41.186 35.234 41.274 ;
        RECT 18.26 41.232 35.188 41.32 ;
        RECT 18.214 41.278 35.142 41.366 ;
        RECT 18.168 41.324 35.096 41.412 ;
        RECT 18.122 41.37 35.05 41.458 ;
        RECT 18.076 41.416 35.004 41.504 ;
        RECT 18.03 41.462 34.958 41.55 ;
        RECT 17.984 41.508 34.912 41.596 ;
        RECT 17.938 41.554 34.866 41.642 ;
        RECT 17.892 41.6 34.82 41.688 ;
        RECT 17.846 41.646 34.774 41.734 ;
        RECT 17.8 41.692 34.728 41.78 ;
        RECT 17.754 41.738 34.682 41.826 ;
        RECT 17.708 41.784 34.636 41.872 ;
        RECT 17.662 41.83 34.59 41.918 ;
        RECT 17.616 41.876 34.544 41.964 ;
        RECT 17.57 41.922 34.498 42.01 ;
        RECT 17.524 41.968 34.452 42.056 ;
        RECT 17.478 42.014 34.406 42.102 ;
        RECT 17.432 42.06 34.36 42.148 ;
        RECT 17.386 42.106 34.314 42.194 ;
        RECT 17.34 42.152 34.268 42.24 ;
        RECT 17.294 42.198 34.222 42.286 ;
        RECT 17.248 42.244 34.176 42.332 ;
        RECT 17.202 42.29 34.13 42.378 ;
        RECT 17.156 42.336 34.084 42.424 ;
        RECT 17.11 42.382 34.038 42.47 ;
        RECT 17.064 42.428 33.992 42.516 ;
        RECT 17.018 42.474 33.946 42.562 ;
        RECT 16.972 42.52 33.9 42.608 ;
        RECT 16.926 42.566 33.854 42.654 ;
        RECT 16.88 42.612 33.808 42.7 ;
        RECT 16.834 42.658 33.762 42.746 ;
        RECT 16.788 42.704 33.716 42.792 ;
        RECT 16.742 42.75 33.67 42.838 ;
        RECT 16.696 42.796 33.624 42.884 ;
        RECT 16.65 42.842 33.578 42.93 ;
        RECT 16.604 42.888 33.532 42.976 ;
        RECT 16.558 42.934 33.486 43.022 ;
        RECT 16.512 42.98 33.44 43.068 ;
        RECT 16.466 43.026 33.394 43.114 ;
        RECT 16.42 43.072 33.348 43.16 ;
        RECT 16.374 43.118 33.302 43.206 ;
        RECT 16.328 43.164 33.256 43.252 ;
        RECT 16.282 43.21 33.21 43.298 ;
        RECT 16.236 43.256 33.164 43.344 ;
        RECT 16.19 43.302 33.118 43.39 ;
        RECT 16.144 43.348 33.072 43.436 ;
        RECT 16.098 43.394 33.026 43.482 ;
        RECT 16.052 43.44 32.98 43.528 ;
        RECT 16.006 43.486 32.934 43.574 ;
        RECT 15.96 43.532 32.888 43.62 ;
        RECT 15.914 43.578 32.842 43.666 ;
        RECT 15.868 43.624 32.796 43.712 ;
        RECT 15.822 43.67 32.75 43.758 ;
        RECT 15.776 43.716 32.704 43.804 ;
        RECT 15.73 43.762 32.658 43.85 ;
        RECT 15.684 43.808 32.612 43.896 ;
        RECT 15.638 43.854 32.566 43.942 ;
        RECT 15.592 43.9 32.52 43.988 ;
        RECT 15.5 43.992 32.474 44.034 ;
        RECT 15.546 43.946 32.474 44.034 ;
        RECT 15.46 44.035 32.428 44.08 ;
        RECT 15.414 44.078 32.382 44.126 ;
        RECT 15.368 44.124 32.336 44.172 ;
        RECT 15.322 44.17 32.29 44.218 ;
        RECT 15.276 44.216 32.244 44.264 ;
        RECT 15.23 44.262 32.198 44.31 ;
        RECT 15.184 44.308 32.152 44.356 ;
        RECT 15.138 44.354 32.106 44.402 ;
        RECT 15.092 44.4 32.06 44.448 ;
        RECT 15.046 44.446 32.014 44.494 ;
        RECT 15 44.492 31.968 44.54 ;
        RECT 14.954 44.538 31.922 44.586 ;
        RECT 14.908 44.584 31.876 44.632 ;
        RECT 14.862 44.63 31.83 44.678 ;
        RECT 14.816 44.676 31.784 44.724 ;
        RECT 14.77 44.722 31.738 44.77 ;
        RECT 14.724 44.768 31.692 44.816 ;
        RECT 14.678 44.814 31.646 44.862 ;
        RECT 14.632 44.86 31.6 44.908 ;
        RECT 14.586 44.906 31.554 44.954 ;
        RECT 14.54 44.952 31.508 45 ;
        RECT 14.494 44.998 31.462 45.046 ;
        RECT 14.448 45.044 31.416 45.092 ;
        RECT 14.402 45.09 31.37 45.138 ;
        RECT 14.356 45.136 31.324 45.184 ;
        RECT 14.31 45.182 31.278 45.23 ;
        RECT 14.264 45.228 31.232 45.276 ;
        RECT 14.218 45.274 31.186 45.322 ;
        RECT 14.172 45.32 31.14 45.368 ;
        RECT 14.126 45.366 31.094 45.414 ;
        RECT 14.08 45.412 31.048 45.46 ;
        RECT 14.034 45.458 31.002 45.506 ;
        RECT 13.988 45.504 30.956 45.552 ;
        RECT 13.942 45.55 30.91 45.598 ;
        RECT 13.896 45.596 30.864 45.644 ;
        RECT 13.85 45.642 30.818 45.69 ;
        RECT 13.804 45.688 30.772 45.736 ;
        RECT 13.758 45.734 30.726 45.782 ;
        RECT 13.712 45.78 30.68 45.828 ;
        RECT 13.666 45.826 30.634 45.874 ;
        RECT 13.62 45.872 30.588 45.92 ;
        RECT 13.574 45.918 30.542 45.966 ;
        RECT 13.528 45.964 30.496 46.012 ;
        RECT 13.482 46.01 30.45 46.058 ;
        RECT 13.436 46.056 30.404 46.104 ;
        RECT 13.39 46.102 30.358 46.15 ;
        RECT 13.344 46.148 30.312 46.196 ;
        RECT 13.298 46.194 30.266 46.242 ;
        RECT 13.252 46.24 30.22 46.288 ;
        RECT 13.206 46.286 30.174 46.334 ;
        RECT 13.16 46.332 30.128 46.38 ;
        RECT 13.114 46.378 30.082 46.426 ;
        RECT 13.068 46.424 30.036 46.472 ;
        RECT 13.022 46.47 29.99 46.518 ;
        RECT 12.976 46.516 29.944 46.564 ;
        RECT 12.93 46.562 29.898 46.61 ;
        RECT 12.884 46.608 29.852 46.656 ;
        RECT 12.838 46.654 29.806 46.702 ;
        RECT 12.792 46.7 29.76 46.748 ;
        RECT 12.746 46.746 29.714 46.794 ;
        RECT 12.7 46.792 29.668 46.84 ;
        RECT 12.654 46.838 29.622 46.886 ;
        RECT 12.608 46.884 29.576 46.932 ;
        RECT 12.562 46.93 29.53 46.978 ;
        RECT 12.516 46.976 29.484 47.024 ;
        RECT 12.47 47.022 29.438 47.07 ;
        RECT 12.424 47.068 29.392 47.116 ;
        RECT 12.378 47.114 29.346 47.162 ;
        RECT 12.332 47.16 29.3 47.208 ;
        RECT 12.286 47.206 29.254 47.254 ;
        RECT 12.24 47.252 29.208 47.3 ;
        RECT 12.194 47.298 29.162 47.346 ;
        RECT 12.148 47.344 29.116 47.392 ;
        RECT 12.102 47.39 29.07 47.438 ;
        RECT 12.056 47.436 29.024 47.484 ;
        RECT 12.01 47.482 28.978 47.53 ;
        RECT 11.964 47.528 28.932 47.576 ;
        RECT 11.918 47.574 28.886 47.622 ;
        RECT 11.872 47.62 28.84 47.668 ;
        RECT 11.826 47.666 28.794 47.714 ;
        RECT 11.78 47.712 28.748 47.76 ;
        RECT 11.734 47.758 28.702 47.806 ;
        RECT 11.688 47.804 28.656 47.852 ;
        RECT 11.642 47.85 28.61 47.898 ;
        RECT 11.596 47.896 28.564 47.944 ;
        RECT 11.55 47.942 28.518 47.99 ;
        RECT 11.504 47.988 28.472 48.036 ;
        RECT 11.458 48.034 28.426 48.082 ;
        RECT 11.412 48.08 28.38 48.128 ;
        RECT 11.366 48.126 28.334 48.174 ;
        RECT 11.32 48.172 28.288 48.22 ;
        RECT 11.274 48.218 28.242 48.266 ;
        RECT 11.228 48.264 28.196 48.312 ;
        RECT 11.182 48.31 28.15 48.358 ;
        RECT 11.136 48.356 28.104 48.404 ;
        RECT 11.09 48.402 28.058 48.45 ;
        RECT 11.044 48.448 28.012 48.496 ;
        RECT 10.998 48.494 27.966 48.542 ;
        RECT 10.952 48.54 27.92 48.588 ;
        RECT 10.906 48.586 27.874 48.634 ;
        RECT 10.86 48.632 27.828 48.68 ;
        RECT 10.814 48.678 27.782 48.726 ;
        RECT 10.768 48.724 27.736 48.772 ;
        RECT 10.722 48.77 27.69 48.818 ;
        RECT 10.676 48.816 27.644 48.864 ;
        RECT 10.63 48.862 27.598 48.91 ;
        RECT 10.584 48.908 27.552 48.956 ;
        RECT 10.538 48.954 27.506 49.002 ;
        RECT 10.492 49 27.46 49.048 ;
        RECT 10.446 49.046 27.414 49.094 ;
        RECT 10.4 49.092 27.368 49.14 ;
        RECT 10.354 49.138 27.322 49.186 ;
        RECT 10.308 49.184 27.276 49.232 ;
        RECT 10.262 49.23 27.23 49.278 ;
        RECT 10.216 49.276 27.184 49.324 ;
        RECT 10.17 49.322 27.138 49.37 ;
        RECT 10.124 49.368 27.092 49.416 ;
        RECT 10.078 49.414 27.046 49.462 ;
    END
  END VSSIO
  OBS
    LAYER MET1 SPACING 0.09 ;
      RECT -20 -20 110 110 ;
    LAYER MET2 SPACING 0.1 ;
      RECT -20 -20 3.325 110 ;
      RECT -20 -20 3.371 55.817 ;
      RECT -20 -20 3.417 55.771 ;
      RECT -20 -20 3.463 55.725 ;
      RECT -20 -20 3.509 55.679 ;
      RECT -20 -20 3.555 55.633 ;
      RECT -20 -20 3.601 55.587 ;
      RECT -20 -20 3.647 55.541 ;
      RECT -20 -20 3.693 55.495 ;
      RECT -20 -20 3.739 55.449 ;
      RECT -20 -20 3.785 55.403 ;
      RECT -20 -20 3.831 55.357 ;
      RECT -20 -20 3.877 55.311 ;
      RECT -20 -20 3.923 55.265 ;
      RECT -20 -20 3.969 55.219 ;
      RECT -20 -20 4.015 55.173 ;
      RECT -20 -20 4.061 55.127 ;
      RECT -20 -20 4.107 55.081 ;
      RECT -20 -20 4.153 55.035 ;
      RECT -20 -20 4.199 54.989 ;
      RECT -20 -20 4.245 54.943 ;
      RECT -20 -20 4.291 54.897 ;
      RECT -20 -20 4.337 54.851 ;
      RECT -20 -20 4.383 54.805 ;
      RECT -20 -20 4.429 54.759 ;
      RECT -20 -20 4.475 54.713 ;
      RECT -20 -20 4.521 54.667 ;
      RECT -20 -20 4.567 54.621 ;
      RECT -20 -20 4.613 54.575 ;
      RECT -20 -20 4.659 54.529 ;
      RECT -20 -20 4.705 54.483 ;
      RECT -20 -20 4.751 54.437 ;
      RECT -20 -20 4.797 54.391 ;
      RECT -20 -20 4.843 54.345 ;
      RECT -20 -20 4.889 54.299 ;
      RECT -20 -20 4.935 54.253 ;
      RECT -20 -20 4.981 54.207 ;
      RECT -20 -20 5.027 54.161 ;
      RECT -20 -20 5.073 54.115 ;
      RECT -20 -20 5.119 54.069 ;
      RECT -20 -20 5.165 54.023 ;
      RECT -20 -20 5.211 53.977 ;
      RECT -20 -20 5.257 53.931 ;
      RECT -20 -20 5.303 53.885 ;
      RECT -20 -20 5.349 53.839 ;
      RECT -20 -20 5.395 53.793 ;
      RECT -20 -20 5.441 53.747 ;
      RECT -20 -20 5.487 53.701 ;
      RECT -20 -20 5.533 53.655 ;
      RECT -20 -20 5.579 53.609 ;
      RECT -20 -20 5.625 53.563 ;
      RECT -20 -20 5.671 53.517 ;
      RECT -20 -20 5.717 53.471 ;
      RECT -20 -20 5.763 53.425 ;
      RECT -20 -20 5.809 53.379 ;
      RECT -20 -20 5.855 53.333 ;
      RECT -20 -20 5.901 53.287 ;
      RECT -20 -20 5.947 53.241 ;
      RECT -20 -20 5.993 53.195 ;
      RECT -20 -20 6.039 53.149 ;
      RECT -20 -20 6.085 53.103 ;
      RECT -20 -20 6.131 53.057 ;
      RECT -20 -20 6.177 53.011 ;
      RECT -20 -20 6.223 52.965 ;
      RECT -20 -20 6.269 52.919 ;
      RECT -20 -20 6.315 52.873 ;
      RECT -20 -20 6.361 52.827 ;
      RECT -20 -20 6.407 52.781 ;
      RECT -20 -20 6.453 52.735 ;
      RECT -20 -20 6.499 52.689 ;
      RECT -20 -20 6.545 52.643 ;
      RECT -20 -20 6.591 52.597 ;
      RECT -20 -20 6.637 52.551 ;
      RECT -20 -20 6.683 52.505 ;
      RECT -20 -20 6.729 52.459 ;
      RECT -20 -20 6.775 52.413 ;
      RECT -20 -20 6.821 52.367 ;
      RECT -20 -20 6.867 52.321 ;
      RECT -20 -20 6.913 52.275 ;
      RECT -20 -20 6.959 52.229 ;
      RECT -20 -20 7.005 52.183 ;
      RECT -20 -20 7.051 52.137 ;
      RECT -20 -20 7.097 52.091 ;
      RECT -20 -20 7.143 52.045 ;
      RECT -20 -20 7.189 51.999 ;
      RECT -20 -20 7.235 51.953 ;
      RECT -20 -20 7.281 51.907 ;
      RECT -20 -20 7.327 51.861 ;
      RECT -20 -20 7.373 51.815 ;
      RECT -20 -20 7.419 51.769 ;
      RECT -20 -20 7.465 51.723 ;
      RECT -20 -20 7.511 51.677 ;
      RECT -20 -20 7.557 51.631 ;
      RECT -20 -20 7.603 51.585 ;
      RECT -20 -20 7.649 51.539 ;
      RECT -20 -20 7.695 51.493 ;
      RECT -20 -20 7.741 51.447 ;
      RECT -20 -20 7.787 51.401 ;
      RECT -20 -20 7.833 51.355 ;
      RECT -20 -20 7.879 51.309 ;
      RECT -20 -20 7.925 51.263 ;
      RECT -20 -20 7.971 51.217 ;
      RECT -20 -20 8.017 51.171 ;
      RECT -20 -20 8.063 51.125 ;
      RECT -20 -20 8.109 51.079 ;
      RECT -20 -20 8.155 51.033 ;
      RECT -20 -20 8.201 50.987 ;
      RECT -20 -20 8.247 50.941 ;
      RECT -20 -20 8.293 50.895 ;
      RECT -20 -20 8.339 50.849 ;
      RECT -20 -20 8.385 50.803 ;
      RECT -20 -20 8.431 50.757 ;
      RECT -20 -20 8.477 50.711 ;
      RECT -20 -20 8.523 50.665 ;
      RECT -20 -20 8.569 50.619 ;
      RECT -20 -20 8.615 50.573 ;
      RECT -20 -20 8.661 50.527 ;
      RECT -20 -20 8.707 50.481 ;
      RECT -20 -20 8.753 50.435 ;
      RECT -20 -20 8.799 50.389 ;
      RECT -20 -20 8.845 50.343 ;
      RECT -20 -20 8.891 50.297 ;
      RECT -20 -20 8.937 50.251 ;
      RECT -20 -20 8.983 50.205 ;
      RECT -20 -20 9.029 50.159 ;
      RECT -20 -20 9.075 50.113 ;
      RECT -20 -20 9.121 50.067 ;
      RECT -20 -20 9.167 50.021 ;
      RECT -20 -20 9.213 49.975 ;
      RECT -20 -20 9.259 49.929 ;
      RECT -20 -20 9.305 49.883 ;
      RECT -20 -20 9.351 49.837 ;
      RECT -20 -20 9.397 49.791 ;
      RECT -20 -20 9.443 49.745 ;
      RECT -20 -20 9.489 49.699 ;
      RECT -20 -20 9.535 49.653 ;
      RECT -20 -20 9.581 49.607 ;
      RECT -20 -20 9.627 49.561 ;
      RECT -20 -20 9.673 49.515 ;
      RECT -20 -20 9.719 49.469 ;
      RECT -20 -20 9.765 49.423 ;
      RECT -20 -20 9.811 49.377 ;
      RECT -20 -20 9.857 49.331 ;
      RECT -20 -20 9.903 49.285 ;
      RECT -20 -20 9.949 49.239 ;
      RECT -20 -20 9.995 49.193 ;
      RECT -20 -20 10.041 49.147 ;
      RECT -20 -20 10.087 49.101 ;
      RECT -20 -20 10.133 49.055 ;
      RECT -20 -20 10.179 49.009 ;
      RECT -20 -20 10.225 48.963 ;
      RECT -20 -20 10.271 48.917 ;
      RECT -20 -20 10.317 48.871 ;
      RECT -20 -20 10.363 48.825 ;
      RECT -20 -20 10.409 48.779 ;
      RECT -20 -20 10.455 48.733 ;
      RECT -20 -20 10.501 48.687 ;
      RECT -20 -20 10.547 48.641 ;
      RECT -20 -20 10.593 48.595 ;
      RECT -20 -20 10.639 48.549 ;
      RECT -20 -20 10.685 48.503 ;
      RECT -20 -20 10.731 48.457 ;
      RECT -20 -20 10.777 48.411 ;
      RECT -20 -20 10.823 48.365 ;
      RECT -20 -20 10.869 48.319 ;
      RECT -20 -20 10.915 48.273 ;
      RECT -20 -20 10.961 48.227 ;
      RECT -20 -20 11.007 48.181 ;
      RECT -20 -20 11.053 48.135 ;
      RECT -20 -20 11.099 48.089 ;
      RECT -20 -20 11.145 48.043 ;
      RECT -20 -20 11.191 47.997 ;
      RECT -20 -20 11.237 47.951 ;
      RECT -20 -20 11.283 47.905 ;
      RECT -20 -20 11.329 47.859 ;
      RECT -20 -20 11.375 47.813 ;
      RECT -20 -20 11.421 47.767 ;
      RECT -20 -20 11.467 47.721 ;
      RECT -20 -20 11.513 47.675 ;
      RECT -20 -20 11.559 47.629 ;
      RECT -20 -20 11.605 47.583 ;
      RECT -20 -20 11.651 47.537 ;
      RECT -20 -20 11.697 47.491 ;
      RECT -20 -20 11.743 47.445 ;
      RECT -20 -20 11.789 47.399 ;
      RECT -20 -20 11.835 47.353 ;
      RECT -20 -20 11.881 47.307 ;
      RECT -20 -20 11.927 47.261 ;
      RECT -20 -20 11.973 47.215 ;
      RECT -20 -20 12.019 47.169 ;
      RECT -20 -20 12.065 47.123 ;
      RECT -20 -20 12.111 47.077 ;
      RECT -20 -20 12.157 47.031 ;
      RECT -20 -20 12.203 46.985 ;
      RECT -20 -20 12.249 46.939 ;
      RECT -20 -20 12.295 46.893 ;
      RECT -20 -20 12.341 46.847 ;
      RECT -20 -20 12.387 46.801 ;
      RECT -20 -20 12.433 46.755 ;
      RECT -20 -20 12.479 46.709 ;
      RECT -20 -20 12.525 46.663 ;
      RECT -20 -20 12.571 46.617 ;
      RECT -20 -20 12.617 46.571 ;
      RECT -20 -20 12.663 46.525 ;
      RECT -20 -20 12.709 46.479 ;
      RECT -20 -20 12.755 46.433 ;
      RECT -20 -20 12.801 46.387 ;
      RECT -20 -20 12.847 46.341 ;
      RECT -20 -20 12.893 46.295 ;
      RECT -20 -20 12.939 46.249 ;
      RECT -20 -20 12.985 46.203 ;
      RECT -20 -20 13.031 46.157 ;
      RECT -20 -20 13.077 46.111 ;
      RECT -20 -20 13.123 46.065 ;
      RECT -20 -20 13.169 46.019 ;
      RECT -20 -20 13.215 45.973 ;
      RECT -20 -20 13.261 45.927 ;
      RECT -20 -20 13.307 45.881 ;
      RECT -20 -20 13.353 45.835 ;
      RECT -20 -20 13.399 45.789 ;
      RECT -20 -20 13.445 45.743 ;
      RECT -20 -20 13.491 45.697 ;
      RECT -20 -20 13.537 45.651 ;
      RECT -20 -20 13.583 45.605 ;
      RECT -20 -20 13.629 45.559 ;
      RECT -20 -20 13.675 45.513 ;
      RECT -20 -20 13.721 45.467 ;
      RECT -20 -20 13.767 45.421 ;
      RECT -20 -20 13.813 45.375 ;
      RECT -20 -20 13.859 45.329 ;
      RECT -20 -20 13.905 45.283 ;
      RECT -20 -20 13.951 45.237 ;
      RECT -20 -20 13.997 45.191 ;
      RECT -20 -20 14.043 45.145 ;
      RECT -20 -20 14.089 45.099 ;
      RECT -20 -20 14.135 45.053 ;
      RECT -20 -20 14.181 45.007 ;
      RECT -20 -20 14.227 44.961 ;
      RECT -20 -20 14.273 44.915 ;
      RECT -20 -20 14.319 44.869 ;
      RECT -20 -20 14.365 44.823 ;
      RECT -20 -20 14.411 44.777 ;
      RECT -20 -20 14.457 44.731 ;
      RECT -20 -20 14.503 44.685 ;
      RECT -20 -20 14.549 44.639 ;
      RECT -20 -20 14.595 44.593 ;
      RECT -20 -20 14.641 44.547 ;
      RECT -20 -20 14.687 44.501 ;
      RECT -20 -20 14.733 44.455 ;
      RECT -20 -20 14.779 44.409 ;
      RECT -20 -20 14.825 44.363 ;
      RECT -20 -20 14.871 44.317 ;
      RECT -20 -20 14.917 44.271 ;
      RECT -20 -20 14.963 44.225 ;
      RECT -20 -20 15.009 44.179 ;
      RECT -20 -20 15.055 44.133 ;
      RECT -20 -20 15.101 44.087 ;
      RECT -20 -20 15.147 44.041 ;
      RECT -20 -20 15.193 43.995 ;
      RECT -20 -20 15.239 43.949 ;
      RECT -20 -20 15.285 43.903 ;
      RECT -20 -20 15.325 43.86 ;
      RECT -20 -20 15.371 43.817 ;
      RECT -20 -20 15.417 43.771 ;
      RECT -20 -20 15.463 43.725 ;
      RECT -20 -20 15.509 43.679 ;
      RECT -20 -20 15.555 43.633 ;
      RECT -20 -20 15.601 43.587 ;
      RECT -20 -20 15.647 43.541 ;
      RECT -20 -20 15.693 43.495 ;
      RECT -20 -20 15.739 43.449 ;
      RECT -20 -20 15.785 43.403 ;
      RECT -20 -20 15.831 43.357 ;
      RECT -20 -20 15.877 43.311 ;
      RECT -20 -20 15.923 43.265 ;
      RECT -20 -20 15.969 43.219 ;
      RECT -20 -20 16.015 43.173 ;
      RECT -20 -20 16.061 43.127 ;
      RECT -20 -20 16.107 43.081 ;
      RECT -20 -20 16.153 43.035 ;
      RECT -20 -20 16.199 42.989 ;
      RECT -20 -20 16.245 42.943 ;
      RECT -20 -20 16.291 42.897 ;
      RECT -20 -20 16.337 42.851 ;
      RECT -20 -20 16.383 42.805 ;
      RECT -20 -20 16.429 42.759 ;
      RECT -20 -20 16.475 42.713 ;
      RECT -20 -20 16.521 42.667 ;
      RECT -20 -20 16.567 42.621 ;
      RECT -20 -20 16.613 42.575 ;
      RECT -20 -20 16.659 42.529 ;
      RECT -20 -20 16.705 42.483 ;
      RECT -20 -20 16.751 42.437 ;
      RECT -20 -20 16.797 42.391 ;
      RECT -20 -20 16.843 42.345 ;
      RECT -20 -20 16.889 42.299 ;
      RECT -20 -20 16.935 42.253 ;
      RECT -20 -20 16.981 42.207 ;
      RECT -20 -20 17.027 42.161 ;
      RECT -20 -20 17.073 42.115 ;
      RECT -20 -20 17.119 42.069 ;
      RECT -20 -20 17.165 42.023 ;
      RECT -20 -20 17.211 41.977 ;
      RECT -20 -20 17.257 41.931 ;
      RECT -20 -20 17.303 41.885 ;
      RECT -20 -20 17.349 41.839 ;
      RECT -20 -20 17.395 41.793 ;
      RECT -20 -20 17.441 41.747 ;
      RECT -20 -20 17.487 41.701 ;
      RECT -20 -20 17.533 41.655 ;
      RECT -20 -20 17.579 41.609 ;
      RECT -20 -20 17.625 41.563 ;
      RECT -20 -20 17.671 41.517 ;
      RECT -20 -20 17.717 41.471 ;
      RECT -20 -20 17.763 41.425 ;
      RECT -20 -20 17.809 41.379 ;
      RECT -20 -20 17.855 41.333 ;
      RECT -20 -20 17.901 41.287 ;
      RECT -20 -20 17.947 41.241 ;
      RECT -20 -20 17.993 41.195 ;
      RECT -20 -20 18.039 41.149 ;
      RECT -20 -20 18.085 41.103 ;
      RECT -20 -20 18.131 41.057 ;
      RECT -20 -20 18.177 41.011 ;
      RECT -20 -20 18.223 40.965 ;
      RECT -20 -20 18.269 40.919 ;
      RECT -20 -20 18.315 40.873 ;
      RECT -20 -20 18.361 40.827 ;
      RECT -20 -20 18.407 40.781 ;
      RECT -20 -20 18.453 40.735 ;
      RECT -20 -20 18.499 40.689 ;
      RECT -20 -20 18.545 40.643 ;
      RECT -20 -20 18.591 40.597 ;
      RECT -20 -20 18.637 40.551 ;
      RECT -20 -20 18.683 40.505 ;
      RECT -20 -20 18.729 40.459 ;
      RECT -20 -20 18.775 40.413 ;
      RECT -20 -20 18.821 40.367 ;
      RECT -20 -20 18.867 40.321 ;
      RECT -20 -20 18.913 40.275 ;
      RECT -20 -20 18.959 40.229 ;
      RECT -20 -20 19.005 40.183 ;
      RECT -20 -20 19.051 40.137 ;
      RECT -20 -20 19.097 40.091 ;
      RECT -20 -20 19.143 40.045 ;
      RECT -20 -20 19.189 39.999 ;
      RECT -20 -20 19.235 39.953 ;
      RECT -20 -20 19.281 39.907 ;
      RECT -20 -20 19.327 39.861 ;
      RECT -20 -20 19.373 39.815 ;
      RECT -20 -20 19.419 39.769 ;
      RECT -20 -20 19.465 39.723 ;
      RECT -20 -20 19.511 39.677 ;
      RECT -20 -20 19.557 39.631 ;
      RECT -20 -20 19.603 39.585 ;
      RECT -20 -20 19.649 39.539 ;
      RECT -20 -20 19.695 39.493 ;
      RECT -20 -20 19.741 39.447 ;
      RECT -20 -20 19.787 39.401 ;
      RECT -20 -20 19.833 39.355 ;
      RECT -20 -20 19.879 39.309 ;
      RECT -20 -20 19.925 39.263 ;
      RECT -20 -20 19.971 39.217 ;
      RECT -20 -20 20.017 39.171 ;
      RECT -20 -20 20.063 39.125 ;
      RECT -20 -20 20.109 39.079 ;
      RECT -20 -20 20.155 39.033 ;
      RECT -20 -20 20.201 38.987 ;
      RECT -20 -20 20.247 38.941 ;
      RECT -20 -20 20.293 38.895 ;
      RECT -20 -20 20.339 38.849 ;
      RECT -20 -20 20.385 38.803 ;
      RECT -20 -20 20.431 38.757 ;
      RECT -20 -20 20.477 38.711 ;
      RECT -20 -20 20.523 38.665 ;
      RECT -20 -20 20.569 38.619 ;
      RECT -20 -20 20.615 38.573 ;
      RECT -20 -20 20.661 38.527 ;
      RECT -20 -20 20.707 38.481 ;
      RECT -20 -20 20.753 38.435 ;
      RECT -20 -20 20.799 38.389 ;
      RECT -20 -20 20.845 38.343 ;
      RECT -20 -20 20.891 38.297 ;
      RECT -20 -20 20.937 38.251 ;
      RECT -20 -20 20.983 38.205 ;
      RECT -20 -20 21.029 38.159 ;
      RECT -20 -20 21.075 38.113 ;
      RECT -20 -20 21.121 38.067 ;
      RECT -20 -20 21.167 38.021 ;
      RECT -20 -20 21.213 37.975 ;
      RECT -20 -20 21.259 37.929 ;
      RECT -20 -20 21.305 37.883 ;
      RECT -20 -20 21.351 37.837 ;
      RECT -20 -20 21.397 37.791 ;
      RECT -20 -20 21.443 37.745 ;
      RECT -20 -20 21.489 37.699 ;
      RECT -20 -20 21.535 37.653 ;
      RECT -20 -20 21.581 37.607 ;
      RECT -20 -20 21.627 37.561 ;
      RECT -20 -20 21.673 37.515 ;
      RECT -20 -20 21.719 37.469 ;
      RECT -20 -20 21.765 37.423 ;
      RECT -20 -20 21.811 37.377 ;
      RECT -20 -20 21.857 37.331 ;
      RECT -20 -20 21.903 37.285 ;
      RECT -20 -20 21.949 37.239 ;
      RECT -20 -20 21.995 37.193 ;
      RECT -20 -20 22.041 37.147 ;
      RECT -20 -20 22.087 37.101 ;
      RECT -20 -20 22.133 37.055 ;
      RECT -20 -20 22.179 37.009 ;
      RECT -20 -20 22.225 36.963 ;
      RECT -20 -20 22.271 36.917 ;
      RECT -20 -20 22.317 36.871 ;
      RECT -20 -20 22.363 36.825 ;
      RECT -20 -20 22.409 36.779 ;
      RECT -20 -20 22.455 36.733 ;
      RECT -20 -20 22.501 36.687 ;
      RECT -20 -20 22.547 36.641 ;
      RECT -20 -20 22.593 36.595 ;
      RECT -20 -20 22.639 36.549 ;
      RECT -20 -20 22.685 36.503 ;
      RECT -20 -20 22.731 36.457 ;
      RECT -20 -20 22.777 36.411 ;
      RECT -20 -20 22.823 36.365 ;
      RECT -20 -20 22.869 36.319 ;
      RECT -20 -20 22.915 36.273 ;
      RECT -20 -20 22.961 36.227 ;
      RECT -20 -20 23.007 36.181 ;
      RECT -20 -20 23.053 36.135 ;
      RECT -20 -20 23.099 36.089 ;
      RECT -20 -20 23.145 36.043 ;
      RECT -20 -20 23.191 35.997 ;
      RECT -20 -20 23.237 35.951 ;
      RECT -20 -20 23.283 35.905 ;
      RECT -20 -20 23.329 35.859 ;
      RECT -20 -20 23.375 35.813 ;
      RECT -20 -20 23.421 35.767 ;
      RECT -20 -20 23.467 35.721 ;
      RECT -20 -20 23.513 35.675 ;
      RECT -20 -20 23.559 35.629 ;
      RECT -20 -20 23.605 35.583 ;
      RECT -20 -20 23.651 35.537 ;
      RECT -20 -20 23.697 35.491 ;
      RECT -20 -20 23.743 35.445 ;
      RECT -20 -20 23.789 35.399 ;
      RECT -20 -20 23.835 35.353 ;
      RECT -20 -20 23.881 35.307 ;
      RECT -20 -20 23.927 35.261 ;
      RECT -20 -20 23.973 35.215 ;
      RECT -20 -20 24.019 35.169 ;
      RECT -20 -20 24.065 35.123 ;
      RECT -20 -20 24.111 35.077 ;
      RECT -20 -20 24.157 35.031 ;
      RECT -20 -20 24.203 34.985 ;
      RECT -20 -20 24.249 34.939 ;
      RECT -20 -20 24.295 34.893 ;
      RECT -20 -20 24.341 34.847 ;
      RECT -20 -20 24.387 34.801 ;
      RECT -20 -20 24.433 34.755 ;
      RECT -20 -20 24.479 34.709 ;
      RECT -20 -20 24.525 34.663 ;
      RECT -20 -20 24.571 34.617 ;
      RECT -20 -20 24.617 34.571 ;
      RECT -20 -20 24.663 34.525 ;
      RECT -20 -20 24.709 34.479 ;
      RECT -20 -20 24.755 34.433 ;
      RECT -20 -20 24.801 34.387 ;
      RECT -20 -20 24.847 34.341 ;
      RECT -20 -20 24.893 34.295 ;
      RECT -20 -20 24.939 34.249 ;
      RECT -20 -20 24.985 34.203 ;
      RECT -20 -20 25.031 34.157 ;
      RECT -20 -20 25.077 34.111 ;
      RECT -20 -20 25.123 34.065 ;
      RECT -20 -20 25.169 34.019 ;
      RECT -20 -20 25.215 33.973 ;
      RECT -20 -20 25.261 33.927 ;
      RECT -20 -20 25.307 33.881 ;
      RECT -20 -20 25.353 33.835 ;
      RECT -20 -20 25.399 33.789 ;
      RECT -20 -20 25.445 33.743 ;
      RECT -20 -20 25.491 33.697 ;
      RECT -20 -20 25.537 33.651 ;
      RECT -20 -20 25.583 33.605 ;
      RECT -20 -20 25.629 33.559 ;
      RECT -20 -20 25.675 33.513 ;
      RECT -20 -20 25.721 33.467 ;
      RECT -20 -20 25.767 33.421 ;
      RECT -20 -20 25.813 33.375 ;
      RECT -20 -20 25.859 33.329 ;
      RECT -20 -20 25.905 33.283 ;
      RECT -20 -20 25.951 33.237 ;
      RECT -20 -20 25.997 33.191 ;
      RECT -20 -20 26.043 33.145 ;
      RECT -20 -20 26.089 33.099 ;
      RECT -20 -20 26.135 33.053 ;
      RECT -20 -20 26.181 33.007 ;
      RECT -20 -20 26.227 32.961 ;
      RECT -20 -20 26.273 32.915 ;
      RECT -20 -20 26.319 32.869 ;
      RECT -20 -20 26.365 32.823 ;
      RECT -20 -20 26.411 32.777 ;
      RECT -20 -20 26.457 32.731 ;
      RECT -20 -20 26.503 32.685 ;
      RECT -20 -20 26.549 32.639 ;
      RECT -20 -20 26.595 32.593 ;
      RECT -20 -20 26.641 32.547 ;
      RECT -20 -20 26.687 32.501 ;
      RECT -20 -20 26.733 32.455 ;
      RECT -20 -20 26.779 32.409 ;
      RECT -20 -20 26.825 32.363 ;
      RECT -20 -20 26.871 32.317 ;
      RECT -20 -20 26.917 32.271 ;
      RECT -20 -20 26.963 32.225 ;
      RECT -20 -20 27.009 32.179 ;
      RECT -20 -20 27.055 32.133 ;
      RECT -20 -20 27.101 32.087 ;
      RECT -20 -20 27.147 32.041 ;
      RECT -20 -20 27.193 31.995 ;
      RECT -20 -20 27.239 31.949 ;
      RECT -20 -20 27.285 31.903 ;
      RECT -20 -20 27.331 31.857 ;
      RECT -20 -20 27.377 31.811 ;
      RECT -20 -20 27.423 31.765 ;
      RECT -20 -20 27.469 31.719 ;
      RECT -20 -20 27.515 31.673 ;
      RECT -20 -20 27.561 31.627 ;
      RECT -20 -20 27.607 31.581 ;
      RECT -20 -20 27.653 31.535 ;
      RECT -20 -20 27.699 31.489 ;
      RECT -20 -20 27.745 31.443 ;
      RECT -20 -20 27.791 31.397 ;
      RECT -20 -20 27.837 31.351 ;
      RECT -20 -20 27.883 31.305 ;
      RECT -20 -20 27.929 31.259 ;
      RECT -20 -20 27.975 31.213 ;
      RECT -20 -20 28.021 31.167 ;
      RECT -20 -20 28.067 31.121 ;
      RECT -20 -20 28.113 31.075 ;
      RECT -20 -20 28.159 31.029 ;
      RECT -20 -20 28.205 30.983 ;
      RECT -20 -20 28.251 30.937 ;
      RECT -20 -20 28.297 30.891 ;
      RECT -20 -20 28.343 30.845 ;
      RECT -20 -20 28.389 30.799 ;
      RECT -20 -20 28.435 30.753 ;
      RECT -20 -20 28.481 30.707 ;
      RECT -20 -20 28.527 30.661 ;
      RECT -20 -20 28.573 30.615 ;
      RECT -20 -20 28.619 30.569 ;
      RECT -20 -20 28.665 30.523 ;
      RECT -20 -20 28.711 30.477 ;
      RECT -20 -20 28.757 30.431 ;
      RECT -20 -20 28.803 30.385 ;
      RECT -20 -20 28.849 30.339 ;
      RECT -20 -20 28.895 30.293 ;
      RECT -20 -20 28.941 30.247 ;
      RECT -20 -20 28.987 30.201 ;
      RECT -20 -20 29.033 30.155 ;
      RECT -20 -20 29.079 30.109 ;
      RECT -20 -20 29.125 30.063 ;
      RECT -20 -20 29.171 30.017 ;
      RECT -20 -20 29.217 29.971 ;
      RECT -20 -20 29.263 29.925 ;
      RECT -20 -20 29.309 29.879 ;
      RECT -20 -20 29.355 29.833 ;
      RECT -20 -20 29.401 29.787 ;
      RECT -20 -20 29.447 29.741 ;
      RECT -20 -20 29.493 29.695 ;
      RECT -20 -20 29.539 29.649 ;
      RECT -20 -20 29.585 29.603 ;
      RECT -20 -20 29.631 29.557 ;
      RECT -20 -20 29.677 29.511 ;
      RECT -20 -20 29.723 29.465 ;
      RECT -20 -20 29.769 29.419 ;
      RECT -20 -20 29.815 29.373 ;
      RECT -20 -20 29.861 29.327 ;
      RECT -20 -20 29.907 29.281 ;
      RECT -20 -20 29.953 29.235 ;
      RECT -20 -20 29.999 29.189 ;
      RECT -20 -20 30.045 29.143 ;
      RECT -20 -20 30.091 29.097 ;
      RECT -20 -20 30.137 29.051 ;
      RECT -20 -20 30.183 29.005 ;
      RECT -20 -20 30.229 28.959 ;
      RECT -20 -20 30.275 28.913 ;
      RECT -20 -20 30.321 28.867 ;
      RECT -20 -20 30.367 28.821 ;
      RECT -20 -20 30.413 28.775 ;
      RECT -20 -20 30.459 28.729 ;
      RECT -20 -20 30.505 28.683 ;
      RECT -20 -20 30.551 28.637 ;
      RECT -20 -20 30.597 28.591 ;
      RECT -20 -20 30.643 28.545 ;
      RECT -20 -20 30.689 28.499 ;
      RECT -20 -20 30.735 28.453 ;
      RECT -20 -20 30.781 28.407 ;
      RECT -20 -20 30.827 28.361 ;
      RECT -20 -20 30.873 28.315 ;
      RECT -20 -20 30.919 28.269 ;
      RECT -20 -20 30.965 28.223 ;
      RECT -20 -20 31.011 28.177 ;
      RECT -20 -20 31.057 28.131 ;
      RECT -20 -20 31.103 28.085 ;
      RECT -20 -20 31.149 28.039 ;
      RECT -20 -20 31.195 27.993 ;
      RECT -20 -20 31.241 27.947 ;
      RECT -20 -20 31.287 27.901 ;
      RECT -20 -20 31.333 27.855 ;
      RECT -20 -20 31.379 27.809 ;
      RECT -20 -20 31.425 27.763 ;
      RECT -20 -20 31.471 27.717 ;
      RECT -20 -20 31.517 27.671 ;
      RECT -20 -20 31.563 27.625 ;
      RECT -20 -20 31.609 27.579 ;
      RECT -20 -20 31.655 27.533 ;
      RECT -20 -20 31.701 27.487 ;
      RECT -20 -20 31.747 27.441 ;
      RECT -20 -20 31.793 27.395 ;
      RECT -20 -20 31.839 27.349 ;
      RECT -20 -20 31.885 27.303 ;
      RECT -20 -20 31.931 27.257 ;
      RECT -20 -20 31.977 27.211 ;
      RECT -20 -20 32.023 27.165 ;
      RECT -20 -20 32.069 27.119 ;
      RECT -20 -20 32.115 27.073 ;
      RECT -20 -20 32.161 27.027 ;
      RECT -20 -20 32.207 26.981 ;
      RECT -20 -20 32.253 26.935 ;
      RECT -20 -20 32.299 26.889 ;
      RECT -20 -20 32.345 26.843 ;
      RECT -20 -20 32.391 26.797 ;
      RECT -20 -20 32.437 26.751 ;
      RECT -20 -20 32.483 26.705 ;
      RECT -20 -20 32.529 26.659 ;
      RECT -20 -20 32.575 26.613 ;
      RECT -20 -20 32.621 26.567 ;
      RECT -20 -20 32.667 26.521 ;
      RECT -20 -20 32.713 26.475 ;
      RECT -20 -20 32.759 26.429 ;
      RECT -20 -20 32.805 26.383 ;
      RECT -20 -20 32.851 26.337 ;
      RECT -20 -20 32.897 26.291 ;
      RECT -20 -20 32.943 26.245 ;
      RECT -20 -20 32.989 26.199 ;
      RECT -20 -20 33.035 26.153 ;
      RECT -20 -20 33.081 26.107 ;
      RECT -20 -20 33.127 26.061 ;
      RECT -20 -20 33.173 26.015 ;
      RECT -20 -20 33.219 25.969 ;
      RECT -20 -20 33.265 25.923 ;
      RECT -20 -20 33.311 25.877 ;
      RECT -20 -20 33.357 25.831 ;
      RECT -20 -20 33.403 25.785 ;
      RECT -20 -20 33.449 25.739 ;
      RECT -20 -20 33.495 25.693 ;
      RECT -20 -20 33.541 25.647 ;
      RECT -20 -20 33.587 25.601 ;
      RECT -20 -20 33.633 25.555 ;
      RECT -20 -20 33.679 25.509 ;
      RECT -20 -20 33.725 25.463 ;
      RECT -20 -20 33.771 25.417 ;
      RECT -20 -20 33.817 25.371 ;
      RECT -20 -20 33.863 25.325 ;
      RECT -20 -20 33.909 25.279 ;
      RECT -20 -20 33.955 25.233 ;
      RECT -20 -20 34.001 25.187 ;
      RECT -20 -20 34.047 25.141 ;
      RECT -20 -20 34.093 25.095 ;
      RECT -20 -20 34.139 25.049 ;
      RECT -20 -20 34.185 25.003 ;
      RECT -20 -20 34.231 24.957 ;
      RECT -20 -20 34.277 24.911 ;
      RECT -20 -20 34.323 24.865 ;
      RECT -20 -20 34.369 24.819 ;
      RECT -20 -20 34.415 24.773 ;
      RECT -20 -20 34.461 24.727 ;
      RECT -20 -20 34.507 24.681 ;
      RECT -20 -20 34.553 24.635 ;
      RECT -20 -20 34.599 24.589 ;
      RECT -20 -20 34.645 24.543 ;
      RECT -20 -20 34.691 24.497 ;
      RECT -20 -20 34.737 24.451 ;
      RECT -20 -20 34.783 24.405 ;
      RECT -20 -20 34.829 24.359 ;
      RECT -20 -20 34.875 24.313 ;
      RECT -20 -20 34.921 24.267 ;
      RECT -20 -20 34.967 24.221 ;
      RECT -20 -20 35.013 24.175 ;
      RECT -20 -20 35.059 24.129 ;
      RECT -20 -20 35.105 24.083 ;
      RECT -20 -20 35.151 24.037 ;
      RECT -20 -20 35.197 23.991 ;
      RECT -20 -20 35.243 23.945 ;
      RECT -20 -20 35.289 23.899 ;
      RECT -20 -20 35.335 23.853 ;
      RECT -20 -20 35.381 23.807 ;
      RECT -20 -20 35.427 23.761 ;
      RECT -20 -20 35.473 23.715 ;
      RECT -20 -20 35.519 23.669 ;
      RECT -20 -20 35.565 23.623 ;
      RECT -20 -20 35.611 23.577 ;
      RECT -20 -20 35.657 23.531 ;
      RECT -20 -20 35.703 23.485 ;
      RECT -20 -20 35.749 23.439 ;
      RECT -20 -20 35.795 23.393 ;
      RECT -20 -20 35.841 23.347 ;
      RECT -20 -20 35.887 23.301 ;
      RECT -20 -20 35.933 23.255 ;
      RECT -20 -20 35.979 23.209 ;
      RECT -20 -20 36.025 23.163 ;
      RECT -20 -20 36.071 23.117 ;
      RECT -20 -20 36.117 23.071 ;
      RECT -20 -20 36.163 23.025 ;
      RECT -20 -20 36.209 22.979 ;
      RECT -20 -20 36.255 22.933 ;
      RECT -20 -20 36.301 22.887 ;
      RECT -20 -20 36.347 22.841 ;
      RECT -20 -20 36.393 22.795 ;
      RECT -20 -20 36.439 22.749 ;
      RECT -20 -20 36.485 22.703 ;
      RECT -20 -20 36.531 22.657 ;
      RECT -20 -20 36.577 22.611 ;
      RECT -20 -20 36.623 22.565 ;
      RECT -20 -20 36.669 22.519 ;
      RECT -20 -20 36.715 22.473 ;
      RECT -20 -20 36.761 22.427 ;
      RECT -20 -20 36.807 22.381 ;
      RECT -20 -20 36.853 22.335 ;
      RECT -20 -20 36.899 22.289 ;
      RECT -20 -20 36.945 22.243 ;
      RECT -20 -20 36.991 22.197 ;
      RECT -20 -20 37.037 22.151 ;
      RECT -20 -20 37.083 22.105 ;
      RECT -20 -20 37.129 22.059 ;
      RECT -20 -20 37.175 22.013 ;
      RECT -20 -20 37.221 21.967 ;
      RECT -20 -20 37.267 21.921 ;
      RECT -20 -20 37.313 21.875 ;
      RECT -20 -20 37.359 21.829 ;
      RECT -20 -20 37.405 21.783 ;
      RECT -20 -20 37.451 21.737 ;
      RECT -20 -20 37.497 21.691 ;
      RECT -20 -20 37.543 21.645 ;
      RECT -20 -20 37.589 21.599 ;
      RECT -20 -20 37.635 21.553 ;
      RECT -20 -20 37.681 21.507 ;
      RECT -20 -20 37.727 21.461 ;
      RECT -20 -20 37.773 21.415 ;
      RECT -20 -20 37.819 21.369 ;
      RECT -20 -20 37.865 21.323 ;
      RECT -20 -20 37.911 21.277 ;
      RECT -20 -20 37.957 21.231 ;
      RECT -20 -20 38.003 21.185 ;
      RECT -20 -20 38.049 21.139 ;
      RECT -20 -20 38.095 21.093 ;
      RECT -20 -20 38.141 21.047 ;
      RECT -20 -20 38.187 21.001 ;
      RECT -20 -20 38.233 20.955 ;
      RECT -20 -20 38.279 20.909 ;
      RECT -20 -20 38.325 20.863 ;
      RECT -20 -20 38.371 20.817 ;
      RECT -20 -20 38.417 20.771 ;
      RECT -20 -20 38.463 20.725 ;
      RECT -20 -20 38.509 20.679 ;
      RECT -20 -20 38.555 20.633 ;
      RECT -20 -20 38.601 20.587 ;
      RECT -20 -20 38.647 20.541 ;
      RECT -20 -20 38.693 20.495 ;
      RECT -20 -20 38.739 20.449 ;
      RECT -20 -20 38.785 20.403 ;
      RECT -20 -20 38.831 20.357 ;
      RECT -20 -20 38.877 20.311 ;
      RECT -20 -20 38.923 20.265 ;
      RECT -20 -20 38.969 20.219 ;
      RECT -20 -20 39.015 20.173 ;
      RECT -20 -20 39.061 20.127 ;
      RECT -20 -20 39.107 20.081 ;
      RECT -20 -20 39.153 20.035 ;
      RECT -20 -20 39.199 19.989 ;
      RECT -20 -20 39.245 19.943 ;
      RECT -20 -20 39.291 19.897 ;
      RECT -20 -20 39.337 19.851 ;
      RECT -20 -20 39.383 19.805 ;
      RECT -20 -20 39.429 19.759 ;
      RECT -20 -20 39.475 19.713 ;
      RECT -20 -20 39.521 19.667 ;
      RECT -20 -20 39.567 19.621 ;
      RECT -20 -20 39.613 19.575 ;
      RECT -20 -20 39.659 19.529 ;
      RECT -20 -20 39.705 19.483 ;
      RECT -20 -20 39.751 19.437 ;
      RECT -20 -20 39.797 19.391 ;
      RECT -20 -20 39.843 19.345 ;
      RECT -20 -20 39.889 19.299 ;
      RECT -20 -20 39.935 19.253 ;
      RECT -20 -20 39.981 19.207 ;
      RECT -20 -20 40.027 19.161 ;
      RECT -20 -20 40.073 19.115 ;
      RECT -20 -20 40.119 19.069 ;
      RECT -20 -20 40.165 19.023 ;
      RECT -20 -20 40.211 18.977 ;
      RECT -20 -20 40.257 18.931 ;
      RECT -20 -20 40.303 18.885 ;
      RECT -20 -20 40.349 18.839 ;
      RECT -20 -20 40.395 18.793 ;
      RECT -20 -20 40.441 18.747 ;
      RECT -20 -20 40.487 18.701 ;
      RECT -20 -20 40.533 18.655 ;
      RECT -20 -20 40.579 18.609 ;
      RECT -20 -20 40.625 18.563 ;
      RECT -20 -20 40.671 18.517 ;
      RECT -20 -20 40.717 18.471 ;
      RECT -20 -20 40.763 18.425 ;
      RECT -20 -20 40.809 18.379 ;
      RECT -20 -20 40.855 18.333 ;
      RECT -20 -20 40.901 18.287 ;
      RECT -20 -20 40.947 18.241 ;
      RECT -20 -20 40.993 18.195 ;
      RECT -20 -20 41.039 18.149 ;
      RECT -20 -20 41.085 18.103 ;
      RECT -20 -20 41.131 18.057 ;
      RECT -20 -20 41.177 18.011 ;
      RECT -20 -20 41.223 17.965 ;
      RECT -20 -20 41.269 17.919 ;
      RECT -20 -20 41.315 17.873 ;
      RECT -20 -20 41.361 17.827 ;
      RECT -20 -20 41.407 17.781 ;
      RECT -20 -20 41.453 17.735 ;
      RECT -20 -20 41.499 17.689 ;
      RECT -20 -20 41.545 17.643 ;
      RECT -20 -20 41.591 17.597 ;
      RECT -20 -20 41.637 17.551 ;
      RECT -20 -20 41.683 17.505 ;
      RECT -20 -20 41.729 17.459 ;
      RECT -20 -20 41.775 17.413 ;
      RECT -20 -20 41.821 17.367 ;
      RECT -20 -20 41.867 17.321 ;
      RECT -20 -20 41.913 17.275 ;
      RECT -20 -20 41.959 17.229 ;
      RECT -20 -20 42.005 17.183 ;
      RECT -20 -20 42.051 17.137 ;
      RECT -20 -20 42.097 17.091 ;
      RECT -20 -20 42.143 17.045 ;
      RECT -20 -20 42.189 16.999 ;
      RECT -20 -20 42.235 16.953 ;
      RECT -20 -20 42.281 16.907 ;
      RECT -20 -20 42.327 16.861 ;
      RECT -20 -20 42.373 16.815 ;
      RECT -20 -20 42.419 16.769 ;
      RECT -20 -20 42.465 16.723 ;
      RECT -20 -20 42.511 16.677 ;
      RECT -20 -20 42.557 16.631 ;
      RECT -20 -20 42.603 16.585 ;
      RECT -20 -20 42.649 16.539 ;
      RECT -20 -20 42.695 16.493 ;
      RECT -20 -20 42.741 16.447 ;
      RECT -20 -20 42.787 16.401 ;
      RECT -20 -20 42.833 16.355 ;
      RECT -20 -20 42.879 16.309 ;
      RECT -20 -20 42.925 16.263 ;
      RECT -20 -20 42.971 16.217 ;
      RECT -20 -20 43.017 16.171 ;
      RECT -20 -20 43.063 16.125 ;
      RECT -20 -20 43.109 16.079 ;
      RECT -20 -20 43.155 16.033 ;
      RECT -20 -20 43.201 15.987 ;
      RECT -20 -20 43.247 15.941 ;
      RECT -20 -20 43.293 15.895 ;
      RECT -20 -20 43.339 15.849 ;
      RECT -20 -20 43.385 15.803 ;
      RECT -20 -20 43.431 15.757 ;
      RECT -20 -20 43.477 15.711 ;
      RECT -20 -20 43.523 15.665 ;
      RECT -20 -20 43.569 15.619 ;
      RECT -20 -20 43.615 15.573 ;
      RECT -20 -20 43.661 15.527 ;
      RECT -20 -20 43.707 15.481 ;
      RECT -20 -20 43.753 15.435 ;
      RECT -20 -20 43.799 15.389 ;
      RECT -20 -20 43.845 15.343 ;
      RECT -20 -20 43.891 15.297 ;
      RECT -20 -20 43.937 15.251 ;
      RECT -20 -20 43.983 15.205 ;
      RECT -20 -20 44.029 15.159 ;
      RECT -20 -20 44.075 15.113 ;
      RECT -20 -20 44.121 15.067 ;
      RECT -20 -20 44.167 15.021 ;
      RECT -20 -20 44.213 14.975 ;
      RECT -20 -20 44.259 14.929 ;
      RECT -20 -20 44.305 14.883 ;
      RECT -20 -20 44.351 14.837 ;
      RECT -20 -20 44.397 14.791 ;
      RECT -20 -20 44.443 14.745 ;
      RECT -20 -20 44.489 14.699 ;
      RECT -20 -20 44.535 14.653 ;
      RECT -20 -20 44.581 14.607 ;
      RECT -20 -20 44.627 14.561 ;
      RECT -20 -20 44.673 14.515 ;
      RECT -20 -20 44.719 14.469 ;
      RECT -20 -20 44.765 14.423 ;
      RECT -20 -20 44.811 14.377 ;
      RECT -20 -20 44.857 14.331 ;
      RECT -20 -20 44.903 14.285 ;
      RECT -20 -20 44.949 14.239 ;
      RECT -20 -20 44.995 14.193 ;
      RECT -20 -20 45.041 14.147 ;
      RECT -20 -20 45.087 14.101 ;
      RECT -20 -20 45.133 14.055 ;
      RECT -20 -20 45.179 14.009 ;
      RECT -20 -20 45.225 13.963 ;
      RECT -20 -20 45.271 13.917 ;
      RECT -20 -20 45.317 13.871 ;
      RECT -20 -20 45.363 13.825 ;
      RECT -20 -20 45.409 13.779 ;
      RECT -20 -20 45.455 13.733 ;
      RECT -20 -20 45.501 13.687 ;
      RECT -20 -20 45.547 13.641 ;
      RECT -20 -20 45.593 13.595 ;
      RECT -20 -20 45.639 13.549 ;
      RECT -20 -20 45.685 13.503 ;
      RECT -20 -20 45.731 13.457 ;
      RECT -20 -20 45.777 13.411 ;
      RECT -20 -20 45.823 13.365 ;
      RECT -20 -20 45.869 13.319 ;
      RECT -20 -20 45.915 13.273 ;
      RECT -20 -20 45.961 13.227 ;
      RECT -20 -20 46.007 13.181 ;
      RECT -20 -20 46.053 13.135 ;
      RECT -20 -20 46.099 13.089 ;
      RECT -20 -20 46.145 13.043 ;
      RECT -20 -20 46.191 12.997 ;
      RECT -20 -20 46.237 12.951 ;
      RECT -20 -20 46.283 12.905 ;
      RECT -20 -20 46.329 12.859 ;
      RECT -20 -20 46.375 12.813 ;
      RECT -20 -20 46.421 12.767 ;
      RECT -20 -20 46.467 12.721 ;
      RECT -20 -20 46.513 12.675 ;
      RECT -20 -20 46.559 12.629 ;
      RECT -20 -20 46.605 12.583 ;
      RECT -20 -20 46.651 12.537 ;
      RECT -20 -20 46.697 12.491 ;
      RECT -20 -20 46.743 12.445 ;
      RECT -20 -20 46.789 12.399 ;
      RECT -20 -20 46.835 12.353 ;
      RECT -20 -20 46.881 12.307 ;
      RECT -20 -20 46.927 12.261 ;
      RECT -20 -20 46.973 12.215 ;
      RECT -20 -20 47.019 12.169 ;
      RECT -20 -20 47.065 12.123 ;
      RECT -20 -20 47.111 12.077 ;
      RECT -20 -20 47.157 12.031 ;
      RECT -20 -20 47.203 11.985 ;
      RECT -20 -20 47.249 11.939 ;
      RECT -20 -20 47.295 11.893 ;
      RECT -20 -20 47.341 11.847 ;
      RECT -20 -20 47.387 11.801 ;
      RECT -20 -20 47.433 11.755 ;
      RECT -20 -20 47.479 11.709 ;
      RECT -20 -20 47.525 11.663 ;
      RECT -20 -20 47.571 11.617 ;
      RECT -20 -20 47.617 11.571 ;
      RECT -20 -20 47.663 11.525 ;
      RECT -20 -20 47.709 11.479 ;
      RECT -20 -20 47.755 11.433 ;
      RECT -20 -20 47.801 11.387 ;
      RECT -20 -20 47.847 11.341 ;
      RECT -20 -20 47.893 11.295 ;
      RECT -20 -20 47.939 11.249 ;
      RECT -20 -20 47.985 11.203 ;
      RECT -20 -20 48.031 11.157 ;
      RECT -20 -20 48.077 11.111 ;
      RECT -20 -20 48.123 11.065 ;
      RECT -20 -20 48.169 11.019 ;
      RECT -20 -20 48.215 10.973 ;
      RECT -20 -20 48.261 10.927 ;
      RECT -20 -20 48.307 10.881 ;
      RECT -20 -20 48.353 10.835 ;
      RECT -20 -20 48.399 10.789 ;
      RECT -20 -20 48.445 10.743 ;
      RECT -20 -20 48.491 10.697 ;
      RECT -20 -20 48.537 10.651 ;
      RECT -20 -20 48.583 10.605 ;
      RECT -20 -20 48.629 10.559 ;
      RECT -20 -20 48.675 10.513 ;
      RECT -20 -20 48.721 10.467 ;
      RECT -20 -20 48.767 10.421 ;
      RECT -20 -20 48.813 10.375 ;
      RECT -20 -20 48.859 10.329 ;
      RECT -20 -20 48.905 10.283 ;
      RECT -20 -20 48.951 10.237 ;
      RECT -20 -20 48.997 10.191 ;
      RECT -20 -20 49.043 10.145 ;
      RECT -20 -20 49.089 10.099 ;
      RECT -20 -20 49.135 10.053 ;
      RECT -20 -20 49.181 10.007 ;
      RECT -20 -20 49.227 9.961 ;
      RECT -20 -20 49.273 9.915 ;
      RECT -20 -20 49.319 9.869 ;
      RECT -20 -20 49.365 9.823 ;
      RECT -20 -20 49.411 9.777 ;
      RECT -20 -20 49.457 9.731 ;
      RECT -20 -20 49.503 9.685 ;
      RECT -20 -20 49.549 9.639 ;
      RECT -20 -20 49.595 9.593 ;
      RECT -20 -20 49.641 9.547 ;
      RECT -20 -20 49.687 9.501 ;
      RECT -20 -20 49.733 9.455 ;
      RECT -20 -20 49.779 9.409 ;
      RECT -20 -20 49.825 9.363 ;
      RECT -20 -20 49.871 9.317 ;
      RECT -20 -20 49.917 9.271 ;
      RECT -20 -20 49.963 9.225 ;
      RECT -20 -20 50.009 9.179 ;
      RECT -20 -20 50.055 9.133 ;
      RECT -20 -20 50.101 9.087 ;
      RECT -20 -20 50.147 9.041 ;
      RECT -20 -20 50.193 8.995 ;
      RECT -20 -20 50.239 8.949 ;
      RECT -20 -20 50.285 8.903 ;
      RECT -20 -20 50.331 8.857 ;
      RECT -20 -20 50.377 8.811 ;
      RECT -20 -20 50.423 8.765 ;
      RECT -20 -20 50.469 8.719 ;
      RECT -20 -20 50.515 8.673 ;
      RECT -20 -20 50.561 8.627 ;
      RECT -20 -20 50.607 8.581 ;
      RECT -20 -20 50.653 8.535 ;
      RECT -20 -20 50.699 8.489 ;
      RECT -20 -20 50.745 8.443 ;
      RECT -20 -20 50.791 8.397 ;
      RECT -20 -20 50.837 8.351 ;
      RECT -20 -20 50.883 8.305 ;
      RECT -20 -20 50.929 8.259 ;
      RECT -20 -20 50.975 8.213 ;
      RECT -20 -20 51.021 8.167 ;
      RECT -20 -20 51.067 8.121 ;
      RECT -20 -20 51.113 8.075 ;
      RECT -20 -20 51.159 8.029 ;
      RECT -20 -20 51.205 7.983 ;
      RECT -20 -20 51.251 7.937 ;
      RECT -20 -20 51.297 7.891 ;
      RECT -20 -20 51.343 7.845 ;
      RECT -20 -20 51.389 7.799 ;
      RECT -20 -20 51.435 7.753 ;
      RECT -20 -20 51.481 7.707 ;
      RECT -20 -20 51.527 7.661 ;
      RECT -20 -20 51.573 7.615 ;
      RECT -20 -20 51.619 7.569 ;
      RECT -20 -20 51.665 7.523 ;
      RECT -20 -20 51.711 7.477 ;
      RECT -20 -20 51.757 7.431 ;
      RECT -20 -20 51.803 7.385 ;
      RECT -20 -20 51.849 7.339 ;
      RECT -20 -20 51.895 7.293 ;
      RECT -20 -20 51.941 7.247 ;
      RECT -20 -20 51.987 7.201 ;
      RECT -20 -20 52.033 7.155 ;
      RECT -20 -20 52.079 7.109 ;
      RECT -20 -20 52.125 7.063 ;
      RECT -20 -20 52.171 7.017 ;
      RECT -20 -20 52.217 6.971 ;
      RECT -20 -20 52.263 6.925 ;
      RECT -20 -20 52.309 6.879 ;
      RECT -20 -20 52.355 6.833 ;
      RECT -20 -20 52.401 6.787 ;
      RECT -20 -20 52.447 6.741 ;
      RECT -20 -20 52.493 6.695 ;
      RECT -20 -20 52.539 6.649 ;
      RECT -20 -20 52.585 6.603 ;
      RECT -20 -20 52.631 6.557 ;
      RECT -20 -20 52.677 6.511 ;
      RECT -20 -20 52.723 6.465 ;
      RECT -20 -20 52.769 6.419 ;
      RECT -20 -20 52.815 6.373 ;
      RECT -20 -20 52.861 6.327 ;
      RECT -20 -20 52.907 6.281 ;
      RECT -20 -20 52.953 6.235 ;
      RECT -20 -20 52.999 6.189 ;
      RECT -20 -20 53.045 6.143 ;
      RECT -20 -20 53.091 6.097 ;
      RECT -20 -20 53.137 6.051 ;
      RECT -20 -20 53.183 6.005 ;
      RECT -20 -20 53.229 5.959 ;
      RECT -20 -20 53.275 5.913 ;
      RECT -20 -20 53.321 5.867 ;
      RECT -20 -20 53.367 5.821 ;
      RECT -20 -20 53.413 5.775 ;
      RECT -20 -20 53.459 5.729 ;
      RECT -20 -20 53.505 5.683 ;
      RECT -20 -20 53.551 5.637 ;
      RECT -20 -20 53.597 5.591 ;
      RECT -20 -20 53.643 5.545 ;
      RECT -20 -20 53.689 5.499 ;
      RECT -20 -20 53.735 5.453 ;
      RECT -20 -20 53.781 5.407 ;
      RECT -20 -20 53.827 5.361 ;
      RECT -20 -20 53.873 5.315 ;
      RECT -20 -20 53.919 5.269 ;
      RECT -20 -20 53.965 5.223 ;
      RECT -20 -20 54.011 5.177 ;
      RECT -20 -20 54.057 5.131 ;
      RECT -20 -20 54.103 5.085 ;
      RECT -20 -20 54.149 5.039 ;
      RECT -20 -20 54.195 4.993 ;
      RECT -20 -20 54.241 4.947 ;
      RECT -20 -20 54.287 4.901 ;
      RECT -20 -20 54.333 4.855 ;
      RECT -20 -20 54.379 4.809 ;
      RECT -20 -20 54.425 4.763 ;
      RECT -20 -20 54.471 4.717 ;
      RECT -20 -20 54.517 4.671 ;
      RECT -20 -20 54.563 4.625 ;
      RECT -20 -20 54.609 4.579 ;
      RECT -20 -20 54.655 4.533 ;
      RECT -20 -20 54.701 4.487 ;
      RECT -20 -20 54.747 4.441 ;
      RECT -20 -20 54.793 4.395 ;
      RECT -20 -20 54.839 4.349 ;
      RECT -20 -20 54.885 4.303 ;
      RECT -20 -20 54.931 4.257 ;
      RECT -20 -20 54.977 4.211 ;
      RECT -20 -20 55.023 4.165 ;
      RECT -20 -20 55.069 4.119 ;
      RECT -20 -20 55.115 4.073 ;
      RECT -20 -20 55.161 4.027 ;
      RECT -20 -20 55.207 3.981 ;
      RECT -20 -20 55.253 3.935 ;
      RECT -20 -20 55.299 3.889 ;
      RECT -20 -20 55.345 3.843 ;
      RECT -20 -20 55.391 3.797 ;
      RECT -20 -20 55.437 3.751 ;
      RECT -20 -20 55.483 3.705 ;
      RECT -20 -20 55.529 3.659 ;
      RECT -20 -20 55.575 3.613 ;
      RECT -20 -20 55.621 3.567 ;
      RECT -20 -20 55.667 3.521 ;
      RECT -20 -20 55.713 3.475 ;
      RECT -20 -20 55.759 3.429 ;
      RECT -20 -20 55.805 3.383 ;
      RECT -20 -20 55.84 3.342 ;
      RECT -20 -20 110 3.325 ;
      RECT 15.675 61.137 16.825 110 ;
      RECT 15.675 61.137 16.871 62.567 ;
      RECT 15.675 61.137 16.917 62.521 ;
      RECT 15.675 61.137 16.963 62.475 ;
      RECT 15.675 61.137 17.009 62.429 ;
      RECT 15.675 61.137 17.055 62.383 ;
      RECT 15.675 61.137 17.101 62.337 ;
      RECT 15.675 61.137 17.147 62.291 ;
      RECT 15.675 61.137 17.193 62.245 ;
      RECT 15.675 61.137 17.239 62.199 ;
      RECT 15.675 61.137 17.285 62.153 ;
      RECT 15.675 61.137 17.331 62.107 ;
      RECT 15.675 61.137 17.377 62.061 ;
      RECT 15.675 61.137 17.423 62.015 ;
      RECT 15.675 61.137 17.469 61.969 ;
      RECT 15.675 61.137 17.515 61.923 ;
      RECT 15.675 61.137 17.561 61.877 ;
      RECT 15.675 61.137 17.607 61.831 ;
      RECT 15.675 61.137 17.653 61.785 ;
      RECT 15.675 61.137 17.699 61.739 ;
      RECT 15.675 61.137 17.745 61.693 ;
      RECT 15.675 61.137 17.791 61.647 ;
      RECT 15.675 61.137 17.837 61.601 ;
      RECT 15.675 61.137 17.883 61.555 ;
      RECT 15.675 61.137 17.929 61.509 ;
      RECT 15.675 61.137 17.975 61.463 ;
      RECT 15.675 61.137 18.021 61.417 ;
      RECT 15.675 61.137 18.067 61.371 ;
      RECT 15.675 61.137 18.113 61.325 ;
      RECT 15.675 61.137 18.159 61.279 ;
      RECT 15.675 61.137 18.205 61.233 ;
      RECT 15.675 61.137 18.251 61.187 ;
      RECT 15.721 61.091 18.297 61.141 ;
      RECT 15.767 61.045 18.343 61.095 ;
      RECT 15.813 60.999 18.389 61.049 ;
      RECT 15.859 60.953 18.435 61.003 ;
      RECT 15.905 60.907 18.481 60.957 ;
      RECT 15.951 60.861 18.527 60.911 ;
      RECT 15.997 60.815 18.573 60.865 ;
      RECT 16.043 60.769 18.619 60.819 ;
      RECT 16.089 60.723 18.665 60.773 ;
      RECT 16.135 60.677 18.711 60.727 ;
      RECT 16.181 60.631 18.757 60.681 ;
      RECT 16.227 60.585 18.803 60.635 ;
      RECT 16.273 60.539 18.849 60.589 ;
      RECT 16.319 60.493 18.895 60.543 ;
      RECT 16.365 60.447 18.941 60.497 ;
      RECT 16.411 60.401 18.987 60.451 ;
      RECT 16.457 60.355 19.033 60.405 ;
      RECT 16.503 60.309 19.079 60.359 ;
      RECT 16.549 60.263 19.125 60.313 ;
      RECT 16.595 60.217 19.171 60.267 ;
      RECT 16.641 60.171 19.217 60.221 ;
      RECT 16.687 60.125 19.263 60.175 ;
      RECT 16.733 60.079 19.309 60.129 ;
      RECT 16.779 60.033 19.355 60.083 ;
      RECT 16.825 59.987 19.401 60.037 ;
      RECT 16.871 59.941 19.447 59.991 ;
      RECT 16.917 59.895 19.493 59.945 ;
      RECT 16.963 59.849 19.539 59.899 ;
      RECT 17.009 59.803 19.585 59.853 ;
      RECT 17.055 59.757 19.631 59.807 ;
      RECT 17.101 59.711 19.677 59.761 ;
      RECT 17.147 59.665 19.723 59.715 ;
      RECT 17.193 59.619 19.769 59.669 ;
      RECT 17.239 59.573 19.815 59.623 ;
      RECT 17.285 59.527 19.861 59.577 ;
      RECT 17.331 59.481 19.907 59.531 ;
      RECT 17.377 59.435 19.953 59.485 ;
      RECT 17.423 59.389 19.999 59.439 ;
      RECT 17.469 59.343 20.045 59.393 ;
      RECT 17.515 59.297 20.091 59.347 ;
      RECT 17.561 59.251 20.137 59.301 ;
      RECT 17.607 59.205 20.183 59.255 ;
      RECT 17.653 59.159 20.229 59.209 ;
      RECT 17.699 59.113 20.275 59.163 ;
      RECT 17.745 59.067 20.321 59.117 ;
      RECT 17.791 59.021 20.367 59.071 ;
      RECT 17.837 58.975 20.413 59.025 ;
      RECT 17.883 58.929 20.459 58.979 ;
      RECT 17.929 58.883 20.505 58.933 ;
      RECT 17.975 58.837 20.551 58.887 ;
      RECT 18.021 58.791 20.597 58.841 ;
      RECT 18.067 58.745 20.643 58.795 ;
      RECT 18.113 58.699 20.689 58.749 ;
      RECT 18.159 58.653 20.735 58.703 ;
      RECT 18.205 58.607 20.781 58.657 ;
      RECT 18.251 58.561 20.827 58.611 ;
      RECT 18.297 58.515 20.873 58.565 ;
      RECT 18.343 58.469 20.919 58.519 ;
      RECT 18.389 58.423 20.965 58.473 ;
      RECT 18.435 58.377 21.011 58.427 ;
      RECT 18.481 58.331 21.057 58.381 ;
      RECT 18.527 58.285 21.103 58.335 ;
      RECT 18.573 58.239 21.149 58.289 ;
      RECT 18.619 58.193 21.195 58.243 ;
      RECT 18.665 58.147 21.241 58.197 ;
      RECT 18.711 58.101 21.287 58.151 ;
      RECT 18.757 58.055 21.333 58.105 ;
      RECT 18.803 58.009 21.379 58.059 ;
      RECT 18.849 57.963 21.425 58.013 ;
      RECT 18.895 57.917 21.471 57.967 ;
      RECT 18.941 57.871 21.517 57.921 ;
      RECT 18.987 57.825 21.563 57.875 ;
      RECT 19.033 57.779 21.609 57.829 ;
      RECT 19.079 57.733 21.655 57.783 ;
      RECT 19.125 57.687 21.701 57.737 ;
      RECT 19.171 57.641 21.747 57.691 ;
      RECT 19.217 57.595 21.793 57.645 ;
      RECT 19.263 57.549 21.839 57.599 ;
      RECT 19.309 57.503 21.885 57.553 ;
      RECT 19.355 57.457 21.931 57.507 ;
      RECT 19.401 57.411 21.977 57.461 ;
      RECT 19.447 57.365 22.023 57.415 ;
      RECT 19.493 57.319 22.069 57.369 ;
      RECT 19.539 57.273 22.115 57.323 ;
      RECT 19.585 57.227 22.161 57.277 ;
      RECT 19.631 57.181 22.207 57.231 ;
      RECT 19.677 57.135 22.253 57.185 ;
      RECT 19.723 57.089 22.299 57.139 ;
      RECT 19.769 57.043 22.345 57.093 ;
      RECT 19.815 56.997 22.391 57.047 ;
      RECT 19.861 56.951 22.437 57.001 ;
      RECT 19.907 56.905 22.483 56.955 ;
      RECT 19.953 56.859 22.529 56.909 ;
      RECT 19.999 56.813 22.575 56.863 ;
      RECT 20.045 56.767 22.621 56.817 ;
      RECT 20.091 56.721 22.667 56.771 ;
      RECT 20.137 56.675 22.713 56.725 ;
      RECT 20.183 56.629 22.759 56.679 ;
      RECT 20.229 56.583 22.805 56.633 ;
      RECT 20.275 56.537 22.851 56.587 ;
      RECT 20.321 56.491 22.897 56.541 ;
      RECT 20.367 56.445 22.943 56.495 ;
      RECT 20.413 56.399 22.989 56.449 ;
      RECT 20.459 56.353 23.035 56.403 ;
      RECT 20.505 56.307 23.081 56.357 ;
      RECT 20.551 56.261 23.127 56.311 ;
      RECT 20.597 56.215 23.173 56.265 ;
      RECT 20.643 56.169 23.219 56.219 ;
      RECT 20.689 56.123 23.265 56.173 ;
      RECT 20.735 56.077 23.311 56.127 ;
      RECT 20.781 56.031 23.357 56.081 ;
      RECT 20.827 55.985 23.403 56.035 ;
      RECT 20.873 55.939 23.449 55.989 ;
      RECT 20.919 55.893 23.495 55.943 ;
      RECT 20.965 55.847 23.541 55.897 ;
      RECT 21.011 55.801 23.587 55.851 ;
      RECT 21.057 55.755 23.633 55.805 ;
      RECT 21.103 55.709 23.679 55.759 ;
      RECT 21.149 55.663 23.725 55.713 ;
      RECT 21.195 55.617 23.771 55.667 ;
      RECT 21.241 55.571 23.817 55.621 ;
      RECT 21.287 55.525 23.863 55.575 ;
      RECT 21.333 55.479 23.909 55.529 ;
      RECT 21.379 55.433 23.955 55.483 ;
      RECT 21.425 55.387 24.001 55.437 ;
      RECT 21.471 55.341 24.047 55.391 ;
      RECT 21.517 55.295 24.093 55.345 ;
      RECT 21.563 55.249 24.139 55.299 ;
      RECT 21.609 55.203 24.185 55.253 ;
      RECT 21.655 55.157 24.231 55.207 ;
      RECT 21.701 55.111 24.277 55.161 ;
      RECT 21.747 55.065 24.323 55.115 ;
      RECT 21.793 55.019 24.369 55.069 ;
      RECT 21.839 54.973 24.415 55.023 ;
      RECT 21.885 54.927 24.461 54.977 ;
      RECT 21.931 54.881 24.507 54.931 ;
      RECT 21.977 54.835 24.553 54.885 ;
      RECT 22.023 54.789 24.599 54.839 ;
      RECT 22.069 54.743 24.645 54.793 ;
      RECT 22.115 54.697 24.691 54.747 ;
      RECT 22.161 54.651 24.737 54.701 ;
      RECT 22.207 54.605 24.783 54.655 ;
      RECT 22.253 54.559 24.829 54.609 ;
      RECT 22.299 54.513 24.875 54.563 ;
      RECT 22.345 54.467 24.921 54.517 ;
      RECT 22.391 54.421 24.967 54.471 ;
      RECT 22.437 54.375 25.013 54.425 ;
      RECT 22.483 54.329 25.059 54.379 ;
      RECT 22.529 54.283 25.105 54.333 ;
      RECT 22.575 54.237 25.151 54.287 ;
      RECT 22.621 54.191 25.197 54.241 ;
      RECT 22.667 54.145 25.243 54.195 ;
      RECT 22.713 54.099 25.289 54.149 ;
      RECT 22.759 54.053 25.335 54.103 ;
      RECT 22.805 54.007 25.381 54.057 ;
      RECT 22.851 53.961 25.427 54.011 ;
      RECT 22.897 53.915 25.473 53.965 ;
      RECT 22.943 53.869 25.519 53.919 ;
      RECT 22.989 53.823 25.565 53.873 ;
      RECT 23.035 53.777 25.611 53.827 ;
      RECT 23.081 53.731 25.657 53.781 ;
      RECT 23.127 53.685 25.703 53.735 ;
      RECT 23.173 53.639 25.749 53.689 ;
      RECT 23.219 53.593 25.795 53.643 ;
      RECT 23.265 53.547 25.841 53.597 ;
      RECT 23.311 53.501 25.887 53.551 ;
      RECT 23.357 53.455 25.933 53.505 ;
      RECT 23.403 53.409 25.979 53.459 ;
      RECT 23.449 53.363 26.025 53.413 ;
      RECT 23.495 53.317 26.071 53.367 ;
      RECT 23.541 53.271 26.117 53.321 ;
      RECT 23.587 53.225 26.163 53.275 ;
      RECT 23.633 53.179 26.209 53.229 ;
      RECT 23.679 53.133 26.255 53.183 ;
      RECT 23.725 53.087 26.301 53.137 ;
      RECT 23.771 53.041 26.347 53.091 ;
      RECT 23.817 52.995 26.393 53.045 ;
      RECT 23.863 52.949 26.439 52.999 ;
      RECT 23.909 52.903 26.485 52.953 ;
      RECT 23.955 52.857 26.531 52.907 ;
      RECT 24.001 52.811 26.577 52.861 ;
      RECT 24.047 52.765 26.623 52.815 ;
      RECT 24.093 52.719 26.669 52.769 ;
      RECT 24.139 52.673 26.715 52.723 ;
      RECT 24.185 52.627 26.761 52.677 ;
      RECT 24.231 52.581 26.807 52.631 ;
      RECT 24.277 52.535 26.853 52.585 ;
      RECT 24.323 52.489 26.899 52.539 ;
      RECT 24.369 52.443 26.945 52.493 ;
      RECT 24.415 52.397 26.991 52.447 ;
      RECT 24.461 52.351 27.037 52.401 ;
      RECT 24.507 52.305 27.083 52.355 ;
      RECT 24.553 52.259 27.129 52.309 ;
      RECT 24.599 52.213 27.175 52.263 ;
      RECT 24.645 52.167 27.221 52.217 ;
      RECT 24.691 52.121 27.267 52.171 ;
      RECT 24.737 52.075 27.313 52.125 ;
      RECT 24.783 52.029 27.359 52.079 ;
      RECT 24.829 51.983 27.405 52.033 ;
      RECT 24.875 51.937 27.451 51.987 ;
      RECT 24.921 51.891 27.497 51.941 ;
      RECT 24.967 51.845 27.543 51.895 ;
      RECT 25.013 51.799 27.589 51.849 ;
      RECT 25.059 51.753 27.635 51.803 ;
      RECT 25.105 51.707 27.681 51.757 ;
      RECT 25.151 51.661 27.727 51.711 ;
      RECT 25.197 51.615 27.773 51.665 ;
      RECT 25.243 51.569 27.819 51.619 ;
      RECT 25.289 51.523 27.865 51.573 ;
      RECT 25.335 51.477 27.911 51.527 ;
      RECT 25.381 51.431 27.957 51.481 ;
      RECT 25.427 51.385 28.003 51.435 ;
      RECT 25.473 51.339 28.049 51.389 ;
      RECT 25.519 51.293 28.095 51.343 ;
      RECT 25.565 51.247 28.141 51.297 ;
      RECT 25.611 51.201 28.187 51.251 ;
      RECT 25.657 51.155 28.233 51.205 ;
      RECT 25.703 51.109 28.279 51.159 ;
      RECT 25.749 51.063 28.325 51.113 ;
      RECT 25.795 51.017 28.371 51.067 ;
      RECT 25.841 50.971 28.417 51.021 ;
      RECT 25.887 50.925 28.463 50.975 ;
      RECT 25.933 50.879 28.509 50.929 ;
      RECT 25.979 50.833 28.555 50.883 ;
      RECT 26.025 50.787 28.601 50.837 ;
      RECT 26.071 50.741 28.647 50.791 ;
      RECT 26.117 50.695 28.693 50.745 ;
      RECT 26.163 50.649 28.739 50.699 ;
      RECT 26.209 50.603 28.785 50.653 ;
      RECT 26.255 50.557 28.825 50.61 ;
      RECT 26.301 50.511 28.871 50.567 ;
      RECT 26.347 50.465 28.917 50.521 ;
      RECT 26.393 50.419 28.963 50.475 ;
      RECT 26.439 50.373 29.009 50.429 ;
      RECT 26.485 50.327 29.055 50.383 ;
      RECT 26.531 50.281 29.101 50.337 ;
      RECT 26.577 50.235 29.147 50.291 ;
      RECT 26.623 50.189 29.193 50.245 ;
      RECT 26.669 50.143 29.239 50.199 ;
      RECT 26.715 50.097 29.285 50.153 ;
      RECT 26.761 50.051 29.331 50.107 ;
      RECT 26.807 50.005 29.377 50.061 ;
      RECT 26.853 49.959 29.423 50.015 ;
      RECT 26.899 49.913 29.469 49.969 ;
      RECT 26.945 49.867 29.515 49.923 ;
      RECT 26.991 49.821 29.561 49.877 ;
      RECT 27.037 49.775 29.607 49.831 ;
      RECT 27.083 49.729 29.653 49.785 ;
      RECT 27.129 49.683 29.699 49.739 ;
      RECT 27.175 49.637 29.745 49.693 ;
      RECT 27.221 49.591 29.791 49.647 ;
      RECT 27.267 49.545 29.837 49.601 ;
      RECT 27.313 49.499 29.883 49.555 ;
      RECT 27.359 49.453 29.929 49.509 ;
      RECT 27.405 49.407 29.975 49.463 ;
      RECT 27.451 49.361 30.021 49.417 ;
      RECT 27.497 49.315 30.067 49.371 ;
      RECT 27.543 49.269 30.113 49.325 ;
      RECT 27.589 49.223 30.159 49.279 ;
      RECT 27.635 49.177 30.205 49.233 ;
      RECT 27.681 49.131 30.251 49.187 ;
      RECT 27.727 49.085 30.297 49.141 ;
      RECT 27.773 49.039 30.343 49.095 ;
      RECT 27.819 48.993 30.389 49.049 ;
      RECT 27.865 48.947 30.435 49.003 ;
      RECT 27.911 48.901 30.481 48.957 ;
      RECT 27.957 48.855 30.527 48.911 ;
      RECT 28.003 48.809 30.573 48.865 ;
      RECT 28.049 48.763 30.619 48.819 ;
      RECT 28.095 48.717 30.665 48.773 ;
      RECT 28.141 48.671 30.711 48.727 ;
      RECT 28.187 48.625 30.757 48.681 ;
      RECT 28.233 48.579 30.803 48.635 ;
      RECT 28.279 48.533 30.849 48.589 ;
      RECT 28.325 48.487 30.895 48.543 ;
      RECT 28.371 48.441 30.941 48.497 ;
      RECT 28.417 48.395 30.987 48.451 ;
      RECT 28.463 48.349 31.033 48.405 ;
      RECT 28.509 48.303 31.079 48.359 ;
      RECT 28.555 48.257 31.125 48.313 ;
      RECT 28.601 48.211 31.171 48.267 ;
      RECT 28.647 48.165 31.217 48.221 ;
      RECT 28.693 48.119 31.263 48.175 ;
      RECT 28.739 48.073 31.309 48.129 ;
      RECT 28.785 48.027 31.355 48.083 ;
      RECT 28.831 47.981 31.401 48.037 ;
      RECT 28.877 47.935 31.447 47.991 ;
      RECT 28.923 47.889 31.493 47.945 ;
      RECT 28.969 47.843 31.539 47.899 ;
      RECT 29.015 47.797 31.585 47.853 ;
      RECT 29.061 47.751 31.631 47.807 ;
      RECT 29.107 47.705 31.677 47.761 ;
      RECT 29.153 47.659 31.723 47.715 ;
      RECT 29.199 47.613 31.769 47.669 ;
      RECT 29.245 47.567 31.815 47.623 ;
      RECT 29.291 47.521 31.861 47.577 ;
      RECT 29.337 47.475 31.907 47.531 ;
      RECT 29.383 47.429 31.953 47.485 ;
      RECT 29.429 47.383 31.999 47.439 ;
      RECT 29.475 47.337 32.045 47.393 ;
      RECT 29.521 47.291 32.091 47.347 ;
      RECT 29.567 47.245 32.137 47.301 ;
      RECT 29.613 47.199 32.183 47.255 ;
      RECT 29.659 47.153 32.229 47.209 ;
      RECT 29.705 47.107 32.275 47.163 ;
      RECT 29.751 47.061 32.321 47.117 ;
      RECT 29.797 47.015 32.367 47.071 ;
      RECT 29.843 46.969 32.413 47.025 ;
      RECT 29.889 46.923 32.459 46.979 ;
      RECT 29.935 46.877 32.505 46.933 ;
      RECT 29.981 46.831 32.551 46.887 ;
      RECT 30.027 46.785 32.597 46.841 ;
      RECT 30.073 46.739 32.643 46.795 ;
      RECT 30.119 46.693 32.689 46.749 ;
      RECT 30.165 46.647 32.735 46.703 ;
      RECT 30.211 46.601 32.781 46.657 ;
      RECT 30.257 46.555 32.827 46.611 ;
      RECT 30.303 46.509 32.873 46.565 ;
      RECT 30.349 46.463 32.919 46.519 ;
      RECT 30.395 46.417 32.965 46.473 ;
      RECT 30.441 46.371 33.011 46.427 ;
      RECT 30.487 46.325 33.057 46.381 ;
      RECT 30.533 46.279 33.103 46.335 ;
      RECT 30.579 46.233 33.149 46.289 ;
      RECT 30.625 46.187 33.195 46.243 ;
      RECT 30.671 46.141 33.241 46.197 ;
      RECT 30.717 46.095 33.287 46.151 ;
      RECT 30.763 46.049 33.333 46.105 ;
      RECT 30.809 46.003 33.379 46.059 ;
      RECT 30.855 45.957 33.425 46.013 ;
      RECT 30.901 45.911 33.471 45.967 ;
      RECT 30.947 45.865 33.517 45.921 ;
      RECT 30.993 45.819 33.563 45.875 ;
      RECT 31.039 45.773 33.609 45.829 ;
      RECT 31.085 45.727 33.655 45.783 ;
      RECT 31.131 45.681 33.701 45.737 ;
      RECT 31.177 45.635 33.747 45.691 ;
      RECT 31.223 45.589 33.793 45.645 ;
      RECT 31.269 45.543 33.839 45.599 ;
      RECT 31.315 45.497 33.885 45.553 ;
      RECT 31.361 45.451 33.931 45.507 ;
      RECT 31.407 45.405 33.977 45.461 ;
      RECT 31.453 45.359 34.023 45.415 ;
      RECT 31.499 45.313 34.069 45.369 ;
      RECT 31.545 45.267 34.115 45.323 ;
      RECT 31.591 45.221 34.161 45.277 ;
      RECT 31.637 45.175 34.207 45.231 ;
      RECT 31.683 45.129 34.253 45.185 ;
      RECT 31.729 45.083 34.299 45.139 ;
      RECT 31.775 45.037 34.345 45.093 ;
      RECT 31.821 44.991 34.391 45.047 ;
      RECT 31.867 44.945 34.437 45.001 ;
      RECT 31.913 44.899 34.483 44.955 ;
      RECT 31.959 44.853 34.529 44.909 ;
      RECT 32.005 44.807 34.575 44.863 ;
      RECT 32.051 44.761 34.621 44.817 ;
      RECT 32.097 44.715 34.667 44.771 ;
      RECT 32.143 44.669 34.713 44.725 ;
      RECT 32.189 44.623 34.759 44.679 ;
      RECT 32.235 44.577 34.805 44.633 ;
      RECT 32.281 44.531 34.851 44.587 ;
      RECT 32.327 44.485 34.897 44.541 ;
      RECT 32.373 44.439 34.943 44.495 ;
      RECT 32.419 44.393 34.989 44.449 ;
      RECT 32.465 44.347 35.035 44.403 ;
      RECT 32.511 44.301 35.081 44.357 ;
      RECT 32.557 44.255 35.127 44.311 ;
      RECT 32.603 44.209 35.173 44.265 ;
      RECT 32.649 44.163 35.219 44.219 ;
      RECT 32.695 44.117 35.265 44.173 ;
      RECT 32.741 44.071 35.311 44.127 ;
      RECT 32.787 44.025 35.357 44.081 ;
      RECT 32.833 43.979 35.403 44.035 ;
      RECT 32.879 43.933 35.449 43.989 ;
      RECT 32.925 43.887 35.495 43.943 ;
      RECT 32.971 43.841 35.541 43.897 ;
      RECT 33.017 43.795 35.587 43.851 ;
      RECT 33.063 43.749 35.633 43.805 ;
      RECT 33.109 43.703 35.679 43.759 ;
      RECT 33.155 43.657 35.725 43.713 ;
      RECT 33.201 43.611 35.771 43.667 ;
      RECT 33.247 43.565 35.817 43.621 ;
      RECT 33.293 43.519 35.863 43.575 ;
      RECT 33.339 43.473 35.909 43.529 ;
      RECT 33.385 43.427 35.955 43.483 ;
      RECT 33.431 43.381 36.001 43.437 ;
      RECT 33.477 43.335 36.047 43.391 ;
      RECT 33.523 43.289 36.093 43.345 ;
      RECT 33.569 43.243 36.139 43.299 ;
      RECT 33.615 43.197 36.185 43.253 ;
      RECT 33.661 43.151 36.231 43.207 ;
      RECT 33.707 43.105 36.277 43.161 ;
      RECT 33.753 43.059 36.323 43.115 ;
      RECT 33.799 43.013 36.369 43.069 ;
      RECT 33.845 42.967 36.415 43.023 ;
      RECT 33.891 42.921 36.461 42.977 ;
      RECT 33.937 42.875 36.507 42.931 ;
      RECT 33.983 42.829 36.553 42.885 ;
      RECT 34.029 42.783 36.599 42.839 ;
      RECT 34.075 42.737 36.645 42.793 ;
      RECT 34.121 42.691 36.691 42.747 ;
      RECT 34.167 42.645 36.737 42.701 ;
      RECT 34.213 42.599 36.783 42.655 ;
      RECT 34.259 42.553 36.829 42.609 ;
      RECT 34.305 42.507 36.875 42.563 ;
      RECT 34.351 42.461 36.921 42.517 ;
      RECT 34.397 42.415 36.967 42.471 ;
      RECT 34.443 42.369 37.013 42.425 ;
      RECT 34.489 42.323 37.059 42.379 ;
      RECT 34.535 42.277 37.105 42.333 ;
      RECT 34.581 42.231 37.151 42.287 ;
      RECT 34.627 42.185 37.197 42.241 ;
      RECT 34.673 42.139 37.243 42.195 ;
      RECT 34.719 42.093 37.289 42.149 ;
      RECT 34.765 42.047 37.335 42.103 ;
      RECT 34.811 42.001 37.381 42.057 ;
      RECT 34.857 41.955 37.427 42.011 ;
      RECT 34.903 41.909 37.473 41.965 ;
      RECT 34.949 41.863 37.519 41.919 ;
      RECT 34.995 41.817 37.565 41.873 ;
      RECT 35.041 41.771 37.611 41.827 ;
      RECT 35.087 41.725 37.657 41.781 ;
      RECT 35.133 41.679 37.703 41.735 ;
      RECT 35.179 41.633 37.749 41.689 ;
      RECT 35.225 41.587 37.795 41.643 ;
      RECT 35.271 41.541 37.841 41.597 ;
      RECT 35.317 41.495 37.887 41.551 ;
      RECT 35.363 41.449 37.933 41.505 ;
      RECT 35.409 41.403 37.979 41.459 ;
      RECT 35.455 41.357 38.025 41.413 ;
      RECT 35.501 41.311 38.071 41.367 ;
      RECT 35.547 41.265 38.117 41.321 ;
      RECT 35.593 41.219 38.163 41.275 ;
      RECT 35.639 41.173 38.209 41.229 ;
      RECT 35.685 41.127 38.255 41.183 ;
      RECT 35.731 41.081 38.301 41.137 ;
      RECT 35.777 41.035 38.347 41.091 ;
      RECT 35.823 40.989 38.393 41.045 ;
      RECT 35.869 40.943 38.439 40.999 ;
      RECT 35.915 40.897 38.485 40.953 ;
      RECT 35.961 40.851 38.531 40.907 ;
      RECT 36.007 40.805 38.577 40.861 ;
      RECT 36.053 40.759 38.623 40.815 ;
      RECT 36.099 40.713 38.669 40.769 ;
      RECT 36.145 40.667 38.715 40.723 ;
      RECT 36.191 40.621 38.761 40.677 ;
      RECT 36.237 40.575 38.807 40.631 ;
      RECT 36.283 40.529 38.853 40.585 ;
      RECT 36.329 40.483 38.899 40.539 ;
      RECT 36.375 40.437 38.945 40.493 ;
      RECT 36.421 40.391 38.991 40.447 ;
      RECT 36.467 40.345 39.037 40.401 ;
      RECT 36.513 40.299 39.083 40.355 ;
      RECT 36.559 40.253 39.129 40.309 ;
      RECT 36.605 40.207 39.175 40.263 ;
      RECT 36.651 40.161 39.221 40.217 ;
      RECT 36.697 40.115 39.267 40.171 ;
      RECT 36.743 40.069 39.313 40.125 ;
      RECT 36.789 40.023 39.359 40.079 ;
      RECT 36.835 39.977 39.405 40.033 ;
      RECT 36.881 39.931 39.451 39.987 ;
      RECT 36.927 39.885 39.497 39.941 ;
      RECT 36.973 39.839 39.543 39.895 ;
      RECT 37.019 39.793 39.589 39.849 ;
      RECT 37.065 39.747 39.635 39.803 ;
      RECT 37.111 39.701 39.681 39.757 ;
      RECT 37.157 39.655 39.727 39.711 ;
      RECT 37.203 39.609 39.773 39.665 ;
      RECT 37.249 39.563 39.819 39.619 ;
      RECT 37.295 39.517 39.865 39.573 ;
      RECT 37.341 39.471 39.911 39.527 ;
      RECT 37.387 39.425 39.957 39.481 ;
      RECT 37.433 39.379 40.003 39.435 ;
      RECT 37.479 39.333 40.049 39.389 ;
      RECT 37.525 39.287 40.095 39.343 ;
      RECT 37.571 39.241 40.141 39.297 ;
      RECT 37.617 39.195 40.187 39.251 ;
      RECT 37.663 39.149 40.233 39.205 ;
      RECT 37.709 39.103 40.279 39.159 ;
      RECT 37.755 39.057 40.325 39.113 ;
      RECT 37.801 39.011 40.371 39.067 ;
      RECT 37.847 38.965 40.417 39.021 ;
      RECT 37.893 38.919 40.463 38.975 ;
      RECT 37.939 38.873 40.509 38.929 ;
      RECT 37.985 38.827 40.555 38.883 ;
      RECT 38.031 38.781 40.601 38.837 ;
      RECT 38.077 38.735 40.647 38.791 ;
      RECT 38.123 38.689 40.693 38.745 ;
      RECT 38.169 38.643 40.739 38.699 ;
      RECT 38.215 38.597 40.785 38.653 ;
      RECT 38.261 38.551 40.831 38.607 ;
      RECT 38.307 38.505 40.877 38.561 ;
      RECT 38.353 38.459 40.923 38.515 ;
      RECT 38.399 38.413 40.969 38.469 ;
      RECT 38.445 38.367 41.015 38.423 ;
      RECT 38.491 38.321 41.061 38.377 ;
      RECT 38.537 38.275 41.107 38.331 ;
      RECT 38.583 38.229 41.153 38.285 ;
      RECT 38.629 38.183 41.199 38.239 ;
      RECT 38.675 38.137 41.245 38.193 ;
      RECT 38.721 38.091 41.291 38.147 ;
      RECT 38.767 38.045 41.337 38.101 ;
      RECT 38.813 37.999 41.383 38.055 ;
      RECT 38.859 37.953 41.429 38.009 ;
      RECT 38.905 37.907 41.475 37.963 ;
      RECT 38.951 37.861 41.521 37.917 ;
      RECT 38.997 37.815 41.567 37.871 ;
      RECT 39.043 37.769 41.613 37.825 ;
      RECT 39.089 37.723 41.659 37.779 ;
      RECT 39.135 37.677 41.705 37.733 ;
      RECT 39.181 37.631 41.751 37.687 ;
      RECT 39.227 37.585 41.797 37.641 ;
      RECT 39.273 37.539 41.843 37.595 ;
      RECT 39.319 37.493 41.889 37.549 ;
      RECT 39.365 37.447 41.935 37.503 ;
      RECT 39.411 37.401 41.981 37.457 ;
      RECT 39.457 37.355 42.027 37.411 ;
      RECT 39.503 37.309 42.073 37.365 ;
      RECT 39.549 37.263 42.119 37.319 ;
      RECT 39.595 37.217 42.165 37.273 ;
      RECT 39.641 37.171 42.211 37.227 ;
      RECT 39.687 37.125 42.257 37.181 ;
      RECT 39.733 37.079 42.303 37.135 ;
      RECT 39.779 37.033 42.349 37.089 ;
      RECT 39.825 36.987 42.395 37.043 ;
      RECT 39.871 36.941 42.441 36.997 ;
      RECT 39.917 36.895 42.487 36.951 ;
      RECT 39.963 36.849 42.533 36.905 ;
      RECT 40.009 36.803 42.579 36.859 ;
      RECT 40.055 36.757 42.625 36.813 ;
      RECT 40.101 36.711 42.671 36.767 ;
      RECT 40.147 36.665 42.717 36.721 ;
      RECT 40.193 36.619 42.763 36.675 ;
      RECT 40.239 36.573 42.809 36.629 ;
      RECT 40.285 36.527 42.855 36.583 ;
      RECT 40.331 36.481 42.901 36.537 ;
      RECT 40.377 36.435 42.947 36.491 ;
      RECT 40.423 36.389 42.993 36.445 ;
      RECT 40.469 36.343 43.039 36.399 ;
      RECT 40.515 36.297 43.085 36.353 ;
      RECT 40.561 36.251 43.131 36.307 ;
      RECT 40.607 36.205 43.177 36.261 ;
      RECT 40.653 36.159 43.223 36.215 ;
      RECT 40.699 36.113 43.269 36.169 ;
      RECT 40.745 36.067 43.315 36.123 ;
      RECT 40.791 36.021 43.361 36.077 ;
      RECT 40.837 35.975 43.407 36.031 ;
      RECT 40.883 35.929 43.453 35.985 ;
      RECT 40.929 35.883 43.499 35.939 ;
      RECT 40.975 35.837 43.545 35.893 ;
      RECT 41.021 35.791 43.591 35.847 ;
      RECT 41.067 35.745 43.637 35.801 ;
      RECT 41.113 35.699 43.683 35.755 ;
      RECT 41.159 35.653 43.729 35.709 ;
      RECT 41.205 35.607 43.775 35.663 ;
      RECT 41.251 35.561 43.821 35.617 ;
      RECT 41.297 35.515 43.867 35.571 ;
      RECT 41.343 35.469 43.913 35.525 ;
      RECT 41.389 35.423 43.959 35.479 ;
      RECT 41.435 35.377 44.005 35.433 ;
      RECT 41.481 35.331 44.051 35.387 ;
      RECT 41.527 35.285 44.097 35.341 ;
      RECT 41.573 35.239 44.143 35.295 ;
      RECT 41.619 35.193 44.189 35.249 ;
      RECT 41.665 35.147 44.235 35.203 ;
      RECT 41.711 35.101 44.281 35.157 ;
      RECT 41.757 35.055 44.327 35.111 ;
      RECT 41.803 35.009 44.373 35.065 ;
      RECT 41.849 34.963 44.419 35.019 ;
      RECT 41.895 34.917 44.465 34.973 ;
      RECT 41.941 34.871 44.511 34.927 ;
      RECT 41.987 34.825 44.557 34.881 ;
      RECT 42.033 34.779 44.603 34.835 ;
      RECT 42.079 34.733 44.649 34.789 ;
      RECT 42.125 34.687 44.695 34.743 ;
      RECT 42.171 34.641 44.741 34.697 ;
      RECT 42.217 34.595 44.787 34.651 ;
      RECT 42.263 34.549 44.833 34.605 ;
      RECT 42.309 34.503 44.879 34.559 ;
      RECT 42.355 34.457 44.925 34.513 ;
      RECT 42.401 34.411 44.971 34.467 ;
      RECT 42.447 34.365 45.017 34.421 ;
      RECT 42.493 34.319 45.063 34.375 ;
      RECT 42.539 34.273 45.109 34.329 ;
      RECT 42.585 34.227 45.155 34.283 ;
      RECT 42.631 34.181 45.201 34.237 ;
      RECT 42.677 34.135 45.247 34.191 ;
      RECT 42.723 34.089 45.293 34.145 ;
      RECT 42.769 34.043 45.339 34.099 ;
      RECT 42.815 33.997 45.385 34.053 ;
      RECT 42.861 33.951 45.431 34.007 ;
      RECT 42.907 33.905 45.477 33.961 ;
      RECT 42.953 33.859 45.523 33.915 ;
      RECT 42.999 33.813 45.569 33.869 ;
      RECT 43.045 33.767 45.615 33.823 ;
      RECT 43.091 33.721 45.661 33.777 ;
      RECT 43.137 33.675 45.707 33.731 ;
      RECT 43.183 33.629 45.753 33.685 ;
      RECT 43.229 33.583 45.799 33.639 ;
      RECT 43.275 33.537 45.845 33.593 ;
      RECT 43.321 33.491 45.891 33.547 ;
      RECT 43.367 33.445 45.937 33.501 ;
      RECT 43.413 33.399 45.983 33.455 ;
      RECT 43.459 33.353 46.029 33.409 ;
      RECT 43.505 33.307 46.075 33.363 ;
      RECT 43.551 33.261 46.121 33.317 ;
      RECT 43.597 33.215 46.167 33.271 ;
      RECT 43.643 33.169 46.213 33.225 ;
      RECT 43.689 33.123 46.259 33.179 ;
      RECT 43.735 33.077 46.305 33.133 ;
      RECT 43.781 33.031 46.351 33.087 ;
      RECT 43.827 32.985 46.397 33.041 ;
      RECT 43.873 32.939 46.443 32.995 ;
      RECT 43.919 32.893 46.489 32.949 ;
      RECT 43.965 32.847 46.535 32.903 ;
      RECT 44.011 32.801 46.581 32.857 ;
      RECT 44.057 32.755 46.627 32.811 ;
      RECT 44.103 32.709 46.673 32.765 ;
      RECT 44.149 32.663 46.719 32.719 ;
      RECT 44.195 32.617 46.765 32.673 ;
      RECT 44.241 32.571 46.811 32.627 ;
      RECT 44.287 32.525 46.857 32.581 ;
      RECT 44.333 32.479 46.903 32.535 ;
      RECT 44.379 32.433 46.949 32.489 ;
      RECT 44.425 32.387 46.995 32.443 ;
      RECT 44.471 32.341 47.041 32.397 ;
      RECT 44.517 32.295 47.087 32.351 ;
      RECT 44.563 32.249 47.133 32.305 ;
      RECT 44.609 32.203 47.179 32.259 ;
      RECT 44.655 32.157 47.225 32.213 ;
      RECT 44.701 32.111 47.271 32.167 ;
      RECT 44.747 32.065 47.317 32.121 ;
      RECT 44.793 32.019 47.363 32.075 ;
      RECT 44.839 31.973 47.409 32.029 ;
      RECT 44.885 31.927 47.455 31.983 ;
      RECT 44.931 31.881 47.501 31.937 ;
      RECT 44.977 31.835 47.547 31.891 ;
      RECT 45.023 31.789 47.593 31.845 ;
      RECT 45.069 31.743 47.639 31.799 ;
      RECT 45.115 31.697 47.685 31.753 ;
      RECT 45.161 31.651 47.731 31.707 ;
      RECT 45.207 31.605 47.777 31.661 ;
      RECT 45.253 31.559 47.823 31.615 ;
      RECT 45.299 31.513 47.869 31.569 ;
      RECT 45.345 31.467 47.915 31.523 ;
      RECT 45.391 31.421 47.961 31.477 ;
      RECT 45.437 31.375 48.007 31.431 ;
      RECT 45.483 31.329 48.053 31.385 ;
      RECT 45.529 31.283 48.099 31.339 ;
      RECT 45.575 31.237 48.145 31.293 ;
      RECT 45.621 31.191 48.191 31.247 ;
      RECT 45.667 31.145 48.237 31.201 ;
      RECT 45.713 31.099 48.283 31.155 ;
      RECT 45.759 31.053 48.329 31.109 ;
      RECT 45.805 31.007 48.375 31.063 ;
      RECT 45.851 30.961 48.421 31.017 ;
      RECT 45.897 30.915 48.467 30.971 ;
      RECT 45.943 30.869 48.513 30.925 ;
      RECT 45.989 30.823 48.559 30.879 ;
      RECT 46.035 30.777 48.605 30.833 ;
      RECT 46.081 30.731 48.651 30.787 ;
      RECT 46.127 30.685 48.697 30.741 ;
      RECT 46.173 30.639 48.743 30.695 ;
      RECT 46.219 30.593 48.789 30.649 ;
      RECT 46.265 30.547 48.835 30.603 ;
      RECT 46.311 30.501 48.881 30.557 ;
      RECT 46.357 30.455 48.927 30.511 ;
      RECT 46.403 30.409 48.973 30.465 ;
      RECT 46.449 30.363 49.019 30.419 ;
      RECT 46.495 30.317 49.065 30.373 ;
      RECT 46.541 30.271 49.111 30.327 ;
      RECT 46.587 30.225 49.157 30.281 ;
      RECT 46.633 30.179 49.203 30.235 ;
      RECT 46.679 30.133 49.249 30.189 ;
      RECT 46.725 30.087 49.295 30.143 ;
      RECT 46.771 30.041 49.341 30.097 ;
      RECT 46.817 29.995 49.387 30.051 ;
      RECT 46.863 29.949 49.433 30.005 ;
      RECT 46.909 29.903 49.479 29.959 ;
      RECT 46.955 29.857 49.525 29.913 ;
      RECT 47.001 29.811 49.571 29.867 ;
      RECT 47.047 29.765 49.617 29.821 ;
      RECT 47.093 29.719 49.663 29.775 ;
      RECT 47.139 29.673 49.709 29.729 ;
      RECT 47.185 29.627 49.755 29.683 ;
      RECT 47.231 29.581 49.801 29.637 ;
      RECT 47.277 29.535 49.847 29.591 ;
      RECT 47.323 29.489 49.893 29.545 ;
      RECT 47.369 29.443 49.939 29.499 ;
      RECT 47.415 29.397 49.985 29.453 ;
      RECT 47.461 29.351 50.031 29.407 ;
      RECT 47.507 29.305 50.077 29.361 ;
      RECT 47.553 29.259 50.123 29.315 ;
      RECT 47.599 29.213 50.169 29.269 ;
      RECT 47.645 29.167 50.215 29.223 ;
      RECT 47.691 29.121 50.261 29.177 ;
      RECT 47.737 29.075 50.307 29.131 ;
      RECT 47.783 29.029 50.353 29.085 ;
      RECT 47.829 28.983 50.399 29.039 ;
      RECT 47.875 28.937 50.445 28.993 ;
      RECT 47.921 28.891 50.491 28.947 ;
      RECT 47.967 28.845 50.537 28.901 ;
      RECT 48.013 28.799 50.583 28.855 ;
      RECT 48.059 28.753 50.629 28.809 ;
      RECT 48.105 28.707 50.675 28.763 ;
      RECT 48.151 28.661 50.721 28.717 ;
      RECT 48.197 28.615 50.767 28.671 ;
      RECT 48.243 28.569 50.813 28.625 ;
      RECT 48.289 28.523 50.859 28.579 ;
      RECT 48.335 28.477 50.905 28.533 ;
      RECT 48.381 28.431 50.951 28.487 ;
      RECT 48.427 28.385 50.997 28.441 ;
      RECT 48.473 28.339 51.043 28.395 ;
      RECT 48.519 28.293 51.089 28.349 ;
      RECT 48.565 28.247 51.135 28.303 ;
      RECT 48.611 28.201 51.181 28.257 ;
      RECT 48.657 28.155 51.227 28.211 ;
      RECT 48.703 28.109 51.273 28.165 ;
      RECT 48.749 28.063 51.319 28.119 ;
      RECT 48.795 28.017 51.365 28.073 ;
      RECT 48.841 27.971 51.411 28.027 ;
      RECT 48.887 27.925 51.457 27.981 ;
      RECT 48.933 27.879 51.503 27.935 ;
      RECT 48.979 27.833 51.549 27.889 ;
      RECT 49.025 27.787 51.595 27.843 ;
      RECT 49.071 27.741 51.641 27.797 ;
      RECT 49.117 27.695 51.687 27.751 ;
      RECT 49.163 27.649 51.733 27.705 ;
      RECT 49.209 27.603 51.779 27.659 ;
      RECT 49.255 27.557 51.825 27.613 ;
      RECT 49.301 27.511 51.871 27.567 ;
      RECT 49.347 27.465 51.917 27.521 ;
      RECT 49.393 27.419 51.963 27.475 ;
      RECT 49.439 27.373 52.009 27.429 ;
      RECT 49.485 27.327 52.055 27.383 ;
      RECT 49.531 27.281 52.101 27.337 ;
      RECT 49.577 27.235 52.147 27.291 ;
      RECT 49.623 27.189 52.193 27.245 ;
      RECT 49.669 27.143 52.239 27.199 ;
      RECT 49.715 27.097 52.285 27.153 ;
      RECT 49.761 27.051 52.331 27.107 ;
      RECT 49.807 27.005 52.377 27.061 ;
      RECT 49.853 26.959 52.423 27.015 ;
      RECT 49.899 26.913 52.469 26.969 ;
      RECT 49.945 26.867 52.515 26.923 ;
      RECT 49.991 26.821 52.561 26.877 ;
      RECT 50.037 26.775 52.607 26.831 ;
      RECT 50.083 26.729 52.653 26.785 ;
      RECT 50.129 26.683 52.699 26.739 ;
      RECT 50.175 26.637 52.745 26.693 ;
      RECT 50.221 26.591 52.791 26.647 ;
      RECT 50.267 26.545 52.837 26.601 ;
      RECT 50.313 26.499 52.883 26.555 ;
      RECT 50.359 26.453 52.929 26.509 ;
      RECT 50.405 26.407 52.975 26.463 ;
      RECT 50.451 26.361 53.021 26.417 ;
      RECT 50.497 26.315 53.067 26.371 ;
      RECT 50.543 26.269 53.113 26.325 ;
      RECT 50.589 26.223 53.159 26.279 ;
      RECT 50.635 26.177 53.205 26.233 ;
      RECT 50.681 26.131 53.251 26.187 ;
      RECT 50.727 26.085 53.297 26.141 ;
      RECT 50.773 26.039 53.343 26.095 ;
      RECT 50.819 25.993 53.389 26.049 ;
      RECT 50.865 25.947 53.435 26.003 ;
      RECT 50.911 25.901 53.481 25.957 ;
      RECT 50.957 25.855 53.527 25.911 ;
      RECT 51.003 25.809 53.573 25.865 ;
      RECT 51.049 25.763 53.619 25.819 ;
      RECT 51.095 25.717 53.665 25.773 ;
      RECT 51.141 25.671 53.711 25.727 ;
      RECT 51.187 25.625 53.757 25.681 ;
      RECT 51.233 25.579 53.803 25.635 ;
      RECT 51.279 25.533 53.849 25.589 ;
      RECT 51.325 25.487 53.895 25.543 ;
      RECT 51.371 25.441 53.941 25.497 ;
      RECT 51.417 25.395 53.987 25.451 ;
      RECT 51.463 25.349 54.033 25.405 ;
      RECT 51.509 25.303 54.079 25.359 ;
      RECT 51.555 25.257 54.125 25.313 ;
      RECT 51.601 25.211 54.171 25.267 ;
      RECT 51.647 25.165 54.217 25.221 ;
      RECT 51.693 25.119 54.263 25.175 ;
      RECT 51.739 25.073 54.309 25.129 ;
      RECT 51.785 25.027 54.355 25.083 ;
      RECT 51.831 24.981 54.401 25.037 ;
      RECT 51.877 24.935 54.447 24.991 ;
      RECT 51.923 24.889 54.493 24.945 ;
      RECT 51.969 24.843 54.539 24.899 ;
      RECT 52.015 24.797 54.585 24.853 ;
      RECT 52.061 24.751 54.631 24.807 ;
      RECT 52.107 24.705 54.677 24.761 ;
      RECT 52.153 24.659 54.723 24.715 ;
      RECT 52.199 24.613 54.769 24.669 ;
      RECT 52.245 24.567 54.815 24.623 ;
      RECT 52.291 24.521 54.861 24.577 ;
      RECT 52.337 24.475 54.907 24.531 ;
      RECT 52.383 24.429 54.953 24.485 ;
      RECT 52.429 24.383 54.999 24.439 ;
      RECT 52.475 24.337 55.045 24.393 ;
      RECT 52.521 24.291 55.091 24.347 ;
      RECT 52.567 24.245 55.137 24.301 ;
      RECT 52.613 24.199 55.183 24.255 ;
      RECT 52.659 24.153 55.229 24.209 ;
      RECT 52.705 24.107 55.275 24.163 ;
      RECT 52.751 24.061 55.321 24.117 ;
      RECT 52.797 24.015 55.367 24.071 ;
      RECT 52.843 23.969 55.413 24.025 ;
      RECT 52.889 23.923 55.459 23.979 ;
      RECT 52.935 23.877 55.505 23.933 ;
      RECT 52.981 23.831 55.551 23.887 ;
      RECT 53.027 23.785 55.597 23.841 ;
      RECT 53.073 23.739 55.643 23.795 ;
      RECT 53.119 23.693 55.689 23.749 ;
      RECT 53.165 23.647 55.735 23.703 ;
      RECT 53.211 23.601 55.781 23.657 ;
      RECT 53.257 23.555 55.827 23.611 ;
      RECT 53.303 23.509 55.873 23.565 ;
      RECT 53.349 23.463 55.919 23.519 ;
      RECT 53.395 23.417 55.965 23.473 ;
      RECT 53.441 23.371 56.011 23.427 ;
      RECT 53.487 23.325 56.057 23.381 ;
      RECT 53.533 23.279 56.103 23.335 ;
      RECT 53.579 23.233 56.149 23.289 ;
      RECT 53.625 23.187 56.195 23.243 ;
      RECT 53.671 23.141 56.241 23.197 ;
      RECT 53.717 23.095 56.287 23.151 ;
      RECT 53.763 23.049 56.333 23.105 ;
      RECT 53.809 23.003 56.379 23.059 ;
      RECT 53.855 22.957 56.425 23.013 ;
      RECT 53.901 22.911 56.471 22.967 ;
      RECT 53.947 22.865 56.517 22.921 ;
      RECT 53.993 22.819 56.563 22.875 ;
      RECT 54.039 22.773 56.609 22.829 ;
      RECT 54.085 22.727 56.655 22.783 ;
      RECT 54.131 22.681 56.701 22.737 ;
      RECT 54.177 22.635 56.747 22.691 ;
      RECT 54.223 22.589 56.793 22.645 ;
      RECT 54.269 22.543 56.839 22.599 ;
      RECT 54.315 22.497 56.885 22.553 ;
      RECT 54.361 22.451 56.931 22.507 ;
      RECT 54.407 22.405 56.977 22.461 ;
      RECT 54.453 22.359 57.023 22.415 ;
      RECT 54.499 22.313 57.069 22.369 ;
      RECT 54.545 22.267 57.115 22.323 ;
      RECT 54.591 22.221 57.161 22.277 ;
      RECT 54.637 22.175 57.207 22.231 ;
      RECT 54.683 22.129 57.253 22.185 ;
      RECT 54.729 22.083 57.299 22.139 ;
      RECT 54.775 22.037 57.345 22.093 ;
      RECT 54.821 21.991 57.391 22.047 ;
      RECT 54.867 21.945 57.437 22.001 ;
      RECT 54.913 21.899 57.483 21.955 ;
      RECT 54.959 21.853 57.529 21.909 ;
      RECT 55.005 21.807 57.575 21.863 ;
      RECT 55.051 21.761 57.621 21.817 ;
      RECT 55.097 21.715 57.667 21.771 ;
      RECT 55.143 21.669 57.713 21.725 ;
      RECT 55.189 21.623 57.759 21.679 ;
      RECT 55.235 21.577 57.805 21.633 ;
      RECT 55.281 21.531 57.851 21.587 ;
      RECT 55.327 21.485 57.897 21.541 ;
      RECT 55.373 21.439 57.943 21.495 ;
      RECT 55.419 21.393 57.989 21.449 ;
      RECT 55.465 21.347 58.035 21.403 ;
      RECT 55.511 21.301 58.081 21.357 ;
      RECT 55.557 21.255 58.127 21.311 ;
      RECT 55.603 21.209 58.173 21.265 ;
      RECT 55.649 21.163 58.219 21.219 ;
      RECT 55.695 21.117 58.265 21.173 ;
      RECT 55.741 21.071 58.311 21.127 ;
      RECT 55.787 21.025 58.357 21.081 ;
      RECT 55.833 20.979 58.403 21.035 ;
      RECT 55.879 20.933 58.449 20.989 ;
      RECT 55.925 20.887 58.495 20.943 ;
      RECT 55.971 20.841 58.541 20.897 ;
      RECT 56.017 20.795 58.587 20.851 ;
      RECT 56.063 20.749 58.633 20.805 ;
      RECT 56.109 20.703 58.679 20.759 ;
      RECT 56.155 20.663 58.725 20.713 ;
      RECT 56.19 20.622 58.771 20.667 ;
      RECT 56.236 20.576 58.817 20.621 ;
      RECT 56.282 20.53 58.863 20.575 ;
      RECT 56.328 20.484 58.909 20.529 ;
      RECT 56.374 20.438 58.955 20.483 ;
      RECT 56.42 20.392 59.001 20.437 ;
      RECT 56.466 20.346 59.047 20.391 ;
      RECT 56.512 20.3 59.093 20.345 ;
      RECT 56.558 20.254 59.139 20.299 ;
      RECT 56.604 20.208 59.185 20.253 ;
      RECT 56.65 20.162 59.231 20.207 ;
      RECT 56.696 20.116 59.277 20.161 ;
      RECT 56.742 20.07 59.323 20.115 ;
      RECT 56.788 20.024 59.369 20.069 ;
      RECT 56.834 19.978 59.415 20.023 ;
      RECT 56.88 19.932 59.461 19.977 ;
      RECT 56.926 19.886 59.507 19.931 ;
      RECT 56.972 19.84 59.553 19.885 ;
      RECT 57.018 19.794 59.599 19.839 ;
      RECT 57.064 19.748 59.645 19.793 ;
      RECT 57.11 19.702 59.691 19.747 ;
      RECT 57.156 19.656 59.737 19.701 ;
      RECT 57.202 19.61 59.783 19.655 ;
      RECT 57.248 19.564 59.829 19.609 ;
      RECT 57.294 19.518 59.875 19.563 ;
      RECT 57.34 19.472 59.921 19.517 ;
      RECT 57.386 19.426 59.967 19.471 ;
      RECT 57.432 19.38 60.013 19.425 ;
      RECT 57.478 19.334 60.059 19.379 ;
      RECT 57.524 19.288 60.105 19.333 ;
      RECT 57.57 19.242 60.151 19.287 ;
      RECT 57.616 19.196 60.197 19.241 ;
      RECT 57.662 19.15 60.243 19.195 ;
      RECT 57.708 19.104 60.289 19.149 ;
      RECT 57.754 19.058 60.335 19.103 ;
      RECT 57.8 19.012 60.381 19.057 ;
      RECT 57.846 18.966 60.427 19.011 ;
      RECT 57.892 18.92 60.473 18.965 ;
      RECT 57.938 18.874 60.519 18.919 ;
      RECT 57.984 18.828 60.565 18.873 ;
      RECT 58.03 18.782 60.611 18.827 ;
      RECT 58.076 18.736 60.657 18.781 ;
      RECT 58.122 18.69 60.703 18.735 ;
      RECT 58.168 18.644 60.749 18.689 ;
      RECT 58.214 18.598 60.795 18.643 ;
      RECT 58.26 18.552 60.841 18.597 ;
      RECT 58.306 18.506 60.887 18.551 ;
      RECT 58.352 18.46 60.933 18.505 ;
      RECT 58.398 18.414 60.979 18.459 ;
      RECT 58.444 18.368 61.025 18.413 ;
      RECT 58.49 18.322 61.071 18.367 ;
      RECT 58.536 18.276 61.117 18.321 ;
      RECT 58.582 18.23 61.163 18.275 ;
      RECT 58.628 18.184 61.209 18.229 ;
      RECT 58.674 18.138 61.255 18.183 ;
      RECT 58.72 18.092 61.301 18.137 ;
      RECT 58.766 18.046 61.347 18.091 ;
      RECT 58.812 18 61.393 18.045 ;
      RECT 58.858 17.954 61.439 17.999 ;
      RECT 58.904 17.908 61.485 17.953 ;
      RECT 58.95 17.862 61.531 17.907 ;
      RECT 58.996 17.816 61.577 17.861 ;
      RECT 59.042 17.77 61.623 17.815 ;
      RECT 59.088 17.724 61.669 17.769 ;
      RECT 59.134 17.678 61.715 17.723 ;
      RECT 59.18 17.632 61.761 17.677 ;
      RECT 59.226 17.586 61.807 17.631 ;
      RECT 59.272 17.54 61.853 17.585 ;
      RECT 59.318 17.494 61.899 17.539 ;
      RECT 59.364 17.448 61.945 17.493 ;
      RECT 59.41 17.402 61.991 17.447 ;
      RECT 59.456 17.356 62.037 17.401 ;
      RECT 59.502 17.31 62.083 17.355 ;
      RECT 59.548 17.264 62.129 17.309 ;
      RECT 59.594 17.218 62.175 17.263 ;
      RECT 59.64 17.172 62.221 17.217 ;
      RECT 59.686 17.126 62.267 17.171 ;
      RECT 59.732 17.08 62.313 17.125 ;
      RECT 59.778 17.034 62.359 17.079 ;
      RECT 59.824 16.988 62.405 17.033 ;
      RECT 59.87 16.942 62.451 16.987 ;
      RECT 59.916 16.896 62.497 16.941 ;
      RECT 59.962 16.85 62.543 16.895 ;
      RECT 60.008 16.804 62.589 16.849 ;
      RECT 61.158 15.675 110 16.825 ;
      RECT 60.054 16.758 110 16.825 ;
      RECT 61.112 15.699 61.163 18.275 ;
      RECT 60.1 16.712 110 16.825 ;
      RECT 61.066 15.746 61.117 18.321 ;
      RECT 60.146 16.666 110 16.825 ;
      RECT 61.02 15.792 61.071 18.367 ;
      RECT 60.192 16.62 110 16.825 ;
      RECT 60.974 15.838 61.025 18.413 ;
      RECT 60.238 16.574 110 16.825 ;
      RECT 60.928 15.884 60.979 18.459 ;
      RECT 60.284 16.528 110 16.825 ;
      RECT 60.882 15.93 60.933 18.505 ;
      RECT 60.33 16.482 110 16.825 ;
      RECT 60.836 15.976 60.887 18.551 ;
      RECT 60.376 16.436 110 16.825 ;
      RECT 60.79 16.022 60.841 18.597 ;
      RECT 60.422 16.39 110 16.825 ;
      RECT 60.744 16.068 60.795 18.643 ;
      RECT 60.468 16.344 110 16.825 ;
      RECT 60.698 16.114 60.749 18.689 ;
      RECT 60.514 16.298 110 16.825 ;
      RECT 60.652 16.16 60.703 18.735 ;
      RECT 60.56 16.252 110 16.825 ;
      RECT 60.606 16.206 60.657 18.781 ;
      RECT 29.175 67.887 30.325 110 ;
      RECT 29.175 67.887 30.371 69.317 ;
      RECT 29.175 67.887 30.417 69.271 ;
      RECT 29.175 67.887 30.463 69.225 ;
      RECT 29.175 67.887 30.509 69.179 ;
      RECT 29.175 67.887 30.555 69.133 ;
      RECT 29.175 67.887 30.601 69.087 ;
      RECT 29.175 67.887 30.647 69.041 ;
      RECT 29.175 67.887 30.693 68.995 ;
      RECT 29.175 67.887 30.739 68.949 ;
      RECT 29.175 67.887 30.785 68.903 ;
      RECT 29.175 67.887 30.831 68.857 ;
      RECT 29.175 67.887 30.877 68.811 ;
      RECT 29.175 67.887 30.923 68.765 ;
      RECT 29.175 67.887 30.969 68.719 ;
      RECT 29.175 67.887 31.015 68.673 ;
      RECT 29.175 67.887 31.061 68.627 ;
      RECT 29.175 67.887 31.107 68.581 ;
      RECT 29.175 67.887 31.153 68.535 ;
      RECT 29.175 67.887 31.199 68.489 ;
      RECT 29.175 67.887 31.245 68.443 ;
      RECT 29.175 67.887 31.291 68.397 ;
      RECT 29.175 67.887 31.337 68.351 ;
      RECT 29.175 67.887 31.383 68.305 ;
      RECT 29.175 67.887 31.429 68.259 ;
      RECT 29.175 67.887 31.475 68.213 ;
      RECT 29.175 67.887 31.521 68.167 ;
      RECT 29.175 67.887 31.567 68.121 ;
      RECT 29.175 67.887 31.613 68.075 ;
      RECT 29.175 67.887 31.659 68.029 ;
      RECT 29.175 67.887 31.705 67.983 ;
      RECT 29.175 67.887 31.751 67.937 ;
      RECT 29.221 67.841 31.797 67.891 ;
      RECT 29.267 67.795 31.843 67.845 ;
      RECT 29.313 67.749 31.889 67.799 ;
      RECT 29.359 67.703 31.935 67.753 ;
      RECT 29.405 67.657 31.981 67.707 ;
      RECT 29.451 67.611 32.027 67.661 ;
      RECT 29.497 67.565 32.073 67.615 ;
      RECT 29.543 67.519 32.119 67.569 ;
      RECT 29.589 67.473 32.165 67.523 ;
      RECT 29.635 67.427 32.211 67.477 ;
      RECT 29.681 67.381 32.257 67.431 ;
      RECT 29.727 67.335 32.303 67.385 ;
      RECT 29.773 67.289 32.349 67.339 ;
      RECT 29.819 67.243 32.395 67.293 ;
      RECT 29.865 67.197 32.441 67.247 ;
      RECT 29.911 67.151 32.487 67.201 ;
      RECT 29.957 67.105 32.533 67.155 ;
      RECT 30.003 67.059 32.579 67.109 ;
      RECT 30.049 67.013 32.625 67.063 ;
      RECT 30.095 66.967 32.671 67.017 ;
      RECT 30.141 66.921 32.717 66.971 ;
      RECT 30.187 66.875 32.763 66.925 ;
      RECT 30.233 66.829 32.809 66.879 ;
      RECT 30.279 66.783 32.855 66.833 ;
      RECT 30.325 66.737 32.901 66.787 ;
      RECT 30.371 66.691 32.947 66.741 ;
      RECT 30.417 66.645 32.993 66.695 ;
      RECT 30.463 66.599 33.039 66.649 ;
      RECT 30.509 66.553 33.085 66.603 ;
      RECT 30.555 66.507 33.131 66.557 ;
      RECT 30.601 66.461 33.177 66.511 ;
      RECT 30.647 66.415 33.223 66.465 ;
      RECT 30.693 66.369 33.269 66.419 ;
      RECT 30.739 66.323 33.315 66.373 ;
      RECT 30.785 66.277 33.361 66.327 ;
      RECT 30.831 66.231 33.407 66.281 ;
      RECT 30.877 66.185 33.453 66.235 ;
      RECT 30.923 66.139 33.499 66.189 ;
      RECT 30.969 66.093 33.545 66.143 ;
      RECT 31.015 66.047 33.591 66.097 ;
      RECT 31.061 66.001 33.637 66.051 ;
      RECT 31.107 65.955 33.683 66.005 ;
      RECT 31.153 65.909 33.729 65.959 ;
      RECT 31.199 65.863 33.775 65.913 ;
      RECT 31.245 65.817 33.821 65.867 ;
      RECT 31.291 65.771 33.867 65.821 ;
      RECT 31.337 65.725 33.913 65.775 ;
      RECT 31.383 65.679 33.959 65.729 ;
      RECT 31.429 65.633 34.005 65.683 ;
      RECT 31.475 65.587 34.051 65.637 ;
      RECT 31.521 65.541 34.097 65.591 ;
      RECT 31.567 65.495 34.143 65.545 ;
      RECT 31.613 65.449 34.189 65.499 ;
      RECT 31.659 65.403 34.235 65.453 ;
      RECT 31.705 65.357 34.281 65.407 ;
      RECT 31.751 65.311 34.327 65.361 ;
      RECT 31.797 65.265 34.373 65.315 ;
      RECT 31.843 65.219 34.419 65.269 ;
      RECT 31.889 65.173 34.465 65.223 ;
      RECT 31.935 65.127 34.511 65.177 ;
      RECT 31.981 65.081 34.557 65.131 ;
      RECT 32.027 65.035 34.603 65.085 ;
      RECT 32.073 64.989 34.649 65.039 ;
      RECT 32.119 64.943 34.695 64.993 ;
      RECT 32.165 64.897 34.741 64.947 ;
      RECT 32.211 64.851 34.787 64.901 ;
      RECT 32.257 64.805 34.833 64.855 ;
      RECT 32.303 64.759 34.879 64.809 ;
      RECT 32.349 64.713 34.925 64.763 ;
      RECT 32.395 64.667 34.971 64.717 ;
      RECT 32.441 64.621 35.017 64.671 ;
      RECT 32.487 64.575 35.063 64.625 ;
      RECT 32.533 64.529 35.109 64.579 ;
      RECT 32.579 64.483 35.155 64.533 ;
      RECT 32.625 64.437 35.201 64.487 ;
      RECT 32.671 64.391 35.247 64.441 ;
      RECT 32.717 64.345 35.293 64.395 ;
      RECT 32.763 64.299 35.339 64.349 ;
      RECT 32.809 64.253 35.385 64.303 ;
      RECT 32.855 64.207 35.431 64.257 ;
      RECT 32.901 64.161 35.477 64.211 ;
      RECT 32.947 64.115 35.523 64.165 ;
      RECT 32.993 64.069 35.569 64.119 ;
      RECT 33.039 64.023 35.615 64.073 ;
      RECT 33.085 63.977 35.661 64.027 ;
      RECT 33.131 63.931 35.707 63.981 ;
      RECT 33.177 63.885 35.753 63.935 ;
      RECT 33.223 63.839 35.799 63.889 ;
      RECT 33.269 63.793 35.845 63.843 ;
      RECT 33.315 63.747 35.891 63.797 ;
      RECT 33.361 63.701 35.937 63.751 ;
      RECT 33.407 63.655 35.983 63.705 ;
      RECT 33.453 63.609 36.029 63.659 ;
      RECT 33.499 63.563 36.075 63.613 ;
      RECT 33.545 63.517 36.121 63.567 ;
      RECT 33.591 63.471 36.167 63.521 ;
      RECT 33.637 63.425 36.213 63.475 ;
      RECT 33.683 63.379 36.259 63.429 ;
      RECT 33.729 63.333 36.305 63.383 ;
      RECT 33.775 63.287 36.351 63.337 ;
      RECT 33.821 63.241 36.397 63.291 ;
      RECT 33.867 63.195 36.443 63.245 ;
      RECT 33.913 63.149 36.489 63.199 ;
      RECT 33.959 63.103 36.535 63.153 ;
      RECT 34.005 63.057 36.581 63.107 ;
      RECT 34.051 63.011 36.627 63.061 ;
      RECT 34.097 62.965 36.673 63.015 ;
      RECT 34.143 62.919 36.719 62.969 ;
      RECT 34.189 62.873 36.765 62.923 ;
      RECT 34.235 62.827 36.811 62.877 ;
      RECT 34.281 62.781 36.857 62.831 ;
      RECT 34.327 62.735 36.903 62.785 ;
      RECT 34.373 62.689 36.949 62.739 ;
      RECT 34.419 62.643 36.995 62.693 ;
      RECT 34.465 62.597 37.041 62.647 ;
      RECT 34.511 62.551 37.087 62.601 ;
      RECT 34.557 62.505 37.133 62.555 ;
      RECT 34.603 62.459 37.179 62.509 ;
      RECT 34.649 62.413 37.225 62.463 ;
      RECT 34.695 62.367 37.271 62.417 ;
      RECT 34.741 62.321 37.317 62.371 ;
      RECT 34.787 62.275 37.363 62.325 ;
      RECT 34.833 62.229 37.409 62.279 ;
      RECT 34.879 62.183 37.455 62.233 ;
      RECT 34.925 62.137 37.501 62.187 ;
      RECT 34.971 62.091 37.547 62.141 ;
      RECT 35.017 62.045 37.593 62.095 ;
      RECT 35.063 61.999 37.639 62.049 ;
      RECT 35.109 61.953 37.685 62.003 ;
      RECT 35.155 61.907 37.731 61.957 ;
      RECT 35.201 61.861 37.777 61.911 ;
      RECT 35.247 61.815 37.823 61.865 ;
      RECT 35.293 61.769 37.869 61.819 ;
      RECT 35.339 61.723 37.915 61.773 ;
      RECT 35.385 61.677 37.961 61.727 ;
      RECT 35.431 61.631 38.007 61.681 ;
      RECT 35.477 61.585 38.053 61.635 ;
      RECT 35.523 61.539 38.099 61.589 ;
      RECT 35.569 61.493 38.145 61.543 ;
      RECT 35.615 61.447 38.191 61.497 ;
      RECT 35.661 61.401 38.237 61.451 ;
      RECT 35.707 61.355 38.283 61.405 ;
      RECT 35.753 61.309 38.329 61.359 ;
      RECT 35.799 61.263 38.375 61.313 ;
      RECT 35.845 61.217 38.421 61.267 ;
      RECT 35.891 61.171 38.467 61.221 ;
      RECT 35.937 61.125 38.513 61.175 ;
      RECT 35.983 61.079 38.559 61.129 ;
      RECT 36.029 61.033 38.605 61.083 ;
      RECT 36.075 60.987 38.651 61.037 ;
      RECT 36.121 60.941 38.697 60.991 ;
      RECT 36.167 60.895 38.743 60.945 ;
      RECT 36.213 60.849 38.789 60.899 ;
      RECT 36.259 60.803 38.835 60.853 ;
      RECT 36.305 60.757 38.881 60.807 ;
      RECT 36.351 60.711 38.927 60.761 ;
      RECT 36.397 60.665 38.973 60.715 ;
      RECT 36.443 60.619 39.019 60.669 ;
      RECT 36.489 60.573 39.065 60.623 ;
      RECT 36.535 60.527 39.111 60.577 ;
      RECT 36.581 60.481 39.157 60.531 ;
      RECT 36.627 60.435 39.203 60.485 ;
      RECT 36.673 60.389 39.249 60.439 ;
      RECT 36.719 60.343 39.295 60.393 ;
      RECT 36.765 60.297 39.341 60.347 ;
      RECT 36.811 60.251 39.387 60.301 ;
      RECT 36.857 60.205 39.433 60.255 ;
      RECT 36.903 60.159 39.479 60.209 ;
      RECT 36.949 60.113 39.525 60.163 ;
      RECT 36.995 60.067 39.571 60.117 ;
      RECT 37.041 60.021 39.617 60.071 ;
      RECT 37.087 59.975 39.663 60.025 ;
      RECT 37.133 59.929 39.709 59.979 ;
      RECT 37.179 59.883 39.755 59.933 ;
      RECT 37.225 59.837 39.801 59.887 ;
      RECT 37.271 59.791 39.847 59.841 ;
      RECT 37.317 59.745 39.893 59.795 ;
      RECT 37.363 59.699 39.939 59.749 ;
      RECT 37.409 59.653 39.985 59.703 ;
      RECT 37.455 59.607 40.031 59.657 ;
      RECT 37.501 59.561 40.077 59.611 ;
      RECT 37.547 59.515 40.123 59.565 ;
      RECT 37.593 59.469 40.169 59.519 ;
      RECT 37.639 59.423 40.215 59.473 ;
      RECT 37.685 59.377 40.261 59.427 ;
      RECT 37.731 59.331 40.307 59.381 ;
      RECT 37.777 59.285 40.353 59.335 ;
      RECT 37.823 59.239 40.399 59.289 ;
      RECT 37.869 59.193 40.445 59.243 ;
      RECT 37.915 59.147 40.491 59.197 ;
      RECT 37.961 59.101 40.537 59.151 ;
      RECT 38.007 59.055 40.583 59.105 ;
      RECT 38.053 59.009 40.629 59.059 ;
      RECT 38.099 58.963 40.675 59.013 ;
      RECT 38.145 58.917 40.721 58.967 ;
      RECT 38.191 58.871 40.767 58.921 ;
      RECT 38.237 58.825 40.813 58.875 ;
      RECT 38.283 58.779 40.859 58.829 ;
      RECT 38.329 58.733 40.905 58.783 ;
      RECT 38.375 58.687 40.951 58.737 ;
      RECT 38.421 58.641 40.997 58.691 ;
      RECT 38.467 58.595 41.043 58.645 ;
      RECT 38.513 58.549 41.089 58.599 ;
      RECT 38.559 58.503 41.135 58.553 ;
      RECT 38.605 58.457 41.181 58.507 ;
      RECT 38.651 58.411 41.227 58.461 ;
      RECT 38.697 58.365 41.273 58.415 ;
      RECT 38.743 58.319 41.319 58.369 ;
      RECT 38.789 58.273 41.365 58.323 ;
      RECT 38.835 58.227 41.411 58.277 ;
      RECT 38.881 58.181 41.457 58.231 ;
      RECT 38.927 58.135 41.503 58.185 ;
      RECT 38.973 58.089 41.549 58.139 ;
      RECT 39.019 58.043 41.595 58.093 ;
      RECT 39.065 57.997 41.641 58.047 ;
      RECT 39.111 57.951 41.687 58.001 ;
      RECT 39.157 57.905 41.733 57.955 ;
      RECT 39.203 57.859 41.779 57.909 ;
      RECT 39.249 57.813 41.825 57.863 ;
      RECT 39.295 57.767 41.871 57.817 ;
      RECT 39.341 57.721 41.917 57.771 ;
      RECT 39.387 57.675 41.963 57.725 ;
      RECT 39.433 57.629 42.009 57.679 ;
      RECT 39.479 57.583 42.055 57.633 ;
      RECT 39.525 57.537 42.101 57.587 ;
      RECT 39.571 57.491 42.147 57.541 ;
      RECT 39.617 57.445 42.193 57.495 ;
      RECT 39.663 57.399 42.239 57.449 ;
      RECT 39.709 57.353 42.285 57.403 ;
      RECT 39.755 57.307 42.325 57.36 ;
      RECT 39.801 57.261 42.371 57.317 ;
      RECT 39.847 57.215 42.417 57.271 ;
      RECT 39.893 57.169 42.463 57.225 ;
      RECT 39.939 57.123 42.509 57.179 ;
      RECT 39.985 57.077 42.555 57.133 ;
      RECT 40.031 57.031 42.601 57.087 ;
      RECT 40.077 56.985 42.647 57.041 ;
      RECT 40.123 56.939 42.693 56.995 ;
      RECT 40.169 56.893 42.739 56.949 ;
      RECT 40.215 56.847 42.785 56.903 ;
      RECT 40.261 56.801 42.831 56.857 ;
      RECT 40.307 56.755 42.877 56.811 ;
      RECT 40.353 56.709 42.923 56.765 ;
      RECT 40.399 56.663 42.969 56.719 ;
      RECT 40.445 56.617 43.015 56.673 ;
      RECT 40.491 56.571 43.061 56.627 ;
      RECT 40.537 56.525 43.107 56.581 ;
      RECT 40.583 56.479 43.153 56.535 ;
      RECT 40.629 56.433 43.199 56.489 ;
      RECT 40.675 56.387 43.245 56.443 ;
      RECT 40.721 56.341 43.291 56.397 ;
      RECT 40.767 56.295 43.337 56.351 ;
      RECT 40.813 56.249 43.383 56.305 ;
      RECT 40.859 56.203 43.429 56.259 ;
      RECT 40.905 56.157 43.475 56.213 ;
      RECT 40.951 56.111 43.521 56.167 ;
      RECT 40.997 56.065 43.567 56.121 ;
      RECT 41.043 56.019 43.613 56.075 ;
      RECT 41.089 55.973 43.659 56.029 ;
      RECT 41.135 55.927 43.705 55.983 ;
      RECT 41.181 55.881 43.751 55.937 ;
      RECT 41.227 55.835 43.797 55.891 ;
      RECT 41.273 55.789 43.843 55.845 ;
      RECT 41.319 55.743 43.889 55.799 ;
      RECT 41.365 55.697 43.935 55.753 ;
      RECT 41.411 55.651 43.981 55.707 ;
      RECT 41.457 55.605 44.027 55.661 ;
      RECT 41.503 55.559 44.073 55.615 ;
      RECT 41.549 55.513 44.119 55.569 ;
      RECT 41.595 55.467 44.165 55.523 ;
      RECT 41.641 55.421 44.211 55.477 ;
      RECT 41.687 55.375 44.257 55.431 ;
      RECT 41.733 55.329 44.303 55.385 ;
      RECT 41.779 55.283 44.349 55.339 ;
      RECT 41.825 55.237 44.395 55.293 ;
      RECT 41.871 55.191 44.441 55.247 ;
      RECT 41.917 55.145 44.487 55.201 ;
      RECT 41.963 55.099 44.533 55.155 ;
      RECT 42.009 55.053 44.579 55.109 ;
      RECT 42.055 55.007 44.625 55.063 ;
      RECT 42.101 54.961 44.671 55.017 ;
      RECT 42.147 54.915 44.717 54.971 ;
      RECT 42.193 54.869 44.763 54.925 ;
      RECT 42.239 54.823 44.809 54.879 ;
      RECT 42.285 54.777 44.855 54.833 ;
      RECT 42.331 54.731 44.901 54.787 ;
      RECT 42.377 54.685 44.947 54.741 ;
      RECT 42.423 54.639 44.993 54.695 ;
      RECT 42.469 54.593 45.039 54.649 ;
      RECT 42.515 54.547 45.085 54.603 ;
      RECT 42.561 54.501 45.131 54.557 ;
      RECT 42.607 54.455 45.177 54.511 ;
      RECT 42.653 54.409 45.223 54.465 ;
      RECT 42.699 54.363 45.269 54.419 ;
      RECT 42.745 54.317 45.315 54.373 ;
      RECT 42.791 54.271 45.361 54.327 ;
      RECT 42.837 54.225 45.407 54.281 ;
      RECT 42.883 54.179 45.453 54.235 ;
      RECT 42.929 54.133 45.499 54.189 ;
      RECT 42.975 54.087 45.545 54.143 ;
      RECT 43.021 54.041 45.591 54.097 ;
      RECT 43.067 53.995 45.637 54.051 ;
      RECT 43.113 53.949 45.683 54.005 ;
      RECT 43.159 53.903 45.729 53.959 ;
      RECT 43.205 53.857 45.775 53.913 ;
      RECT 43.251 53.811 45.821 53.867 ;
      RECT 43.297 53.765 45.867 53.821 ;
      RECT 43.343 53.719 45.913 53.775 ;
      RECT 43.389 53.673 45.959 53.729 ;
      RECT 43.435 53.627 46.005 53.683 ;
      RECT 43.481 53.581 46.051 53.637 ;
      RECT 43.527 53.535 46.097 53.591 ;
      RECT 43.573 53.489 46.143 53.545 ;
      RECT 43.619 53.443 46.189 53.499 ;
      RECT 43.665 53.397 46.235 53.453 ;
      RECT 43.711 53.351 46.281 53.407 ;
      RECT 43.757 53.305 46.327 53.361 ;
      RECT 43.803 53.259 46.373 53.315 ;
      RECT 43.849 53.213 46.419 53.269 ;
      RECT 43.895 53.167 46.465 53.223 ;
      RECT 43.941 53.121 46.511 53.177 ;
      RECT 43.987 53.075 46.557 53.131 ;
      RECT 44.033 53.029 46.603 53.085 ;
      RECT 44.079 52.983 46.649 53.039 ;
      RECT 44.125 52.937 46.695 52.993 ;
      RECT 44.171 52.891 46.741 52.947 ;
      RECT 44.217 52.845 46.787 52.901 ;
      RECT 44.263 52.799 46.833 52.855 ;
      RECT 44.309 52.753 46.879 52.809 ;
      RECT 44.355 52.707 46.925 52.763 ;
      RECT 44.401 52.661 46.971 52.717 ;
      RECT 44.447 52.615 47.017 52.671 ;
      RECT 44.493 52.569 47.063 52.625 ;
      RECT 44.539 52.523 47.109 52.579 ;
      RECT 44.585 52.477 47.155 52.533 ;
      RECT 44.631 52.431 47.201 52.487 ;
      RECT 44.677 52.385 47.247 52.441 ;
      RECT 44.723 52.339 47.293 52.395 ;
      RECT 44.769 52.293 47.339 52.349 ;
      RECT 44.815 52.247 47.385 52.303 ;
      RECT 44.861 52.201 47.431 52.257 ;
      RECT 44.907 52.155 47.477 52.211 ;
      RECT 44.953 52.109 47.523 52.165 ;
      RECT 44.999 52.063 47.569 52.119 ;
      RECT 45.045 52.017 47.615 52.073 ;
      RECT 45.091 51.971 47.661 52.027 ;
      RECT 45.137 51.925 47.707 51.981 ;
      RECT 45.183 51.879 47.753 51.935 ;
      RECT 45.229 51.833 47.799 51.889 ;
      RECT 45.275 51.787 47.845 51.843 ;
      RECT 45.321 51.741 47.891 51.797 ;
      RECT 45.367 51.695 47.937 51.751 ;
      RECT 45.413 51.649 47.983 51.705 ;
      RECT 45.459 51.603 48.029 51.659 ;
      RECT 45.505 51.557 48.075 51.613 ;
      RECT 45.551 51.511 48.121 51.567 ;
      RECT 45.597 51.465 48.167 51.521 ;
      RECT 45.643 51.419 48.213 51.475 ;
      RECT 45.689 51.373 48.259 51.429 ;
      RECT 45.735 51.327 48.305 51.383 ;
      RECT 45.781 51.281 48.351 51.337 ;
      RECT 45.827 51.235 48.397 51.291 ;
      RECT 45.873 51.189 48.443 51.245 ;
      RECT 45.919 51.143 48.489 51.199 ;
      RECT 45.965 51.097 48.535 51.153 ;
      RECT 46.011 51.051 48.581 51.107 ;
      RECT 46.057 51.005 48.627 51.061 ;
      RECT 46.103 50.959 48.673 51.015 ;
      RECT 46.149 50.913 48.719 50.969 ;
      RECT 46.195 50.867 48.765 50.923 ;
      RECT 46.241 50.821 48.811 50.877 ;
      RECT 46.287 50.775 48.857 50.831 ;
      RECT 46.333 50.729 48.903 50.785 ;
      RECT 46.379 50.683 48.949 50.739 ;
      RECT 46.425 50.637 48.995 50.693 ;
      RECT 46.471 50.591 49.041 50.647 ;
      RECT 46.517 50.545 49.087 50.601 ;
      RECT 46.563 50.499 49.133 50.555 ;
      RECT 46.609 50.453 49.179 50.509 ;
      RECT 46.655 50.407 49.225 50.463 ;
      RECT 46.701 50.361 49.271 50.417 ;
      RECT 46.747 50.315 49.317 50.371 ;
      RECT 46.793 50.269 49.363 50.325 ;
      RECT 46.839 50.223 49.409 50.279 ;
      RECT 46.885 50.177 49.455 50.233 ;
      RECT 46.931 50.131 49.501 50.187 ;
      RECT 46.977 50.085 49.547 50.141 ;
      RECT 47.023 50.039 49.593 50.095 ;
      RECT 47.069 49.993 49.639 50.049 ;
      RECT 47.115 49.947 49.685 50.003 ;
      RECT 47.161 49.901 49.731 49.957 ;
      RECT 47.207 49.855 49.777 49.911 ;
      RECT 47.253 49.809 49.823 49.865 ;
      RECT 47.299 49.763 49.869 49.819 ;
      RECT 47.345 49.717 49.915 49.773 ;
      RECT 47.391 49.671 49.961 49.727 ;
      RECT 47.437 49.625 50.007 49.681 ;
      RECT 47.483 49.579 50.053 49.635 ;
      RECT 47.529 49.533 50.099 49.589 ;
      RECT 47.575 49.487 50.145 49.543 ;
      RECT 47.621 49.441 50.191 49.497 ;
      RECT 47.667 49.395 50.237 49.451 ;
      RECT 47.713 49.349 50.283 49.405 ;
      RECT 47.759 49.303 50.329 49.359 ;
      RECT 47.805 49.257 50.375 49.313 ;
      RECT 47.851 49.211 50.421 49.267 ;
      RECT 47.897 49.165 50.467 49.221 ;
      RECT 47.943 49.119 50.513 49.175 ;
      RECT 47.989 49.073 50.559 49.129 ;
      RECT 48.035 49.027 50.605 49.083 ;
      RECT 48.081 48.981 50.651 49.037 ;
      RECT 48.127 48.935 50.697 48.991 ;
      RECT 48.173 48.889 50.743 48.945 ;
      RECT 48.219 48.843 50.789 48.899 ;
      RECT 48.265 48.797 50.835 48.853 ;
      RECT 48.311 48.751 50.881 48.807 ;
      RECT 48.357 48.705 50.927 48.761 ;
      RECT 48.403 48.659 50.973 48.715 ;
      RECT 48.449 48.613 51.019 48.669 ;
      RECT 48.495 48.567 51.065 48.623 ;
      RECT 48.541 48.521 51.111 48.577 ;
      RECT 48.587 48.475 51.157 48.531 ;
      RECT 48.633 48.429 51.203 48.485 ;
      RECT 48.679 48.383 51.249 48.439 ;
      RECT 48.725 48.337 51.295 48.393 ;
      RECT 48.771 48.291 51.341 48.347 ;
      RECT 48.817 48.245 51.387 48.301 ;
      RECT 48.863 48.199 51.433 48.255 ;
      RECT 48.909 48.153 51.479 48.209 ;
      RECT 48.955 48.107 51.525 48.163 ;
      RECT 49.001 48.061 51.571 48.117 ;
      RECT 49.047 48.015 51.617 48.071 ;
      RECT 49.093 47.969 51.663 48.025 ;
      RECT 49.139 47.923 51.709 47.979 ;
      RECT 49.185 47.877 51.755 47.933 ;
      RECT 49.231 47.831 51.801 47.887 ;
      RECT 49.277 47.785 51.847 47.841 ;
      RECT 49.323 47.739 51.893 47.795 ;
      RECT 49.369 47.693 51.939 47.749 ;
      RECT 49.415 47.647 51.985 47.703 ;
      RECT 49.461 47.601 52.031 47.657 ;
      RECT 49.507 47.555 52.077 47.611 ;
      RECT 49.553 47.509 52.123 47.565 ;
      RECT 49.599 47.463 52.169 47.519 ;
      RECT 49.645 47.417 52.215 47.473 ;
      RECT 49.691 47.371 52.261 47.427 ;
      RECT 49.737 47.325 52.307 47.381 ;
      RECT 49.783 47.279 52.353 47.335 ;
      RECT 49.829 47.233 52.399 47.289 ;
      RECT 49.875 47.187 52.445 47.243 ;
      RECT 49.921 47.141 52.491 47.197 ;
      RECT 49.967 47.095 52.537 47.151 ;
      RECT 50.013 47.049 52.583 47.105 ;
      RECT 50.059 47.003 52.629 47.059 ;
      RECT 50.105 46.957 52.675 47.013 ;
      RECT 50.151 46.911 52.721 46.967 ;
      RECT 50.197 46.865 52.767 46.921 ;
      RECT 50.243 46.819 52.813 46.875 ;
      RECT 50.289 46.773 52.859 46.829 ;
      RECT 50.335 46.727 52.905 46.783 ;
      RECT 50.381 46.681 52.951 46.737 ;
      RECT 50.427 46.635 52.997 46.691 ;
      RECT 50.473 46.589 53.043 46.645 ;
      RECT 50.519 46.543 53.089 46.599 ;
      RECT 50.565 46.497 53.135 46.553 ;
      RECT 50.611 46.451 53.181 46.507 ;
      RECT 50.657 46.405 53.227 46.461 ;
      RECT 50.703 46.359 53.273 46.415 ;
      RECT 50.749 46.313 53.319 46.369 ;
      RECT 50.795 46.267 53.365 46.323 ;
      RECT 50.841 46.221 53.411 46.277 ;
      RECT 50.887 46.175 53.457 46.231 ;
      RECT 50.933 46.129 53.503 46.185 ;
      RECT 50.979 46.083 53.549 46.139 ;
      RECT 51.025 46.037 53.595 46.093 ;
      RECT 51.071 45.991 53.641 46.047 ;
      RECT 51.117 45.945 53.687 46.001 ;
      RECT 51.163 45.899 53.733 45.955 ;
      RECT 51.209 45.853 53.779 45.909 ;
      RECT 51.255 45.807 53.825 45.863 ;
      RECT 51.301 45.761 53.871 45.817 ;
      RECT 51.347 45.715 53.917 45.771 ;
      RECT 51.393 45.669 53.963 45.725 ;
      RECT 51.439 45.623 54.009 45.679 ;
      RECT 51.485 45.577 54.055 45.633 ;
      RECT 51.531 45.531 54.101 45.587 ;
      RECT 51.577 45.485 54.147 45.541 ;
      RECT 51.623 45.439 54.193 45.495 ;
      RECT 51.669 45.393 54.239 45.449 ;
      RECT 51.715 45.347 54.285 45.403 ;
      RECT 51.761 45.301 54.331 45.357 ;
      RECT 51.807 45.255 54.377 45.311 ;
      RECT 51.853 45.209 54.423 45.265 ;
      RECT 51.899 45.163 54.469 45.219 ;
      RECT 51.945 45.117 54.515 45.173 ;
      RECT 51.991 45.071 54.561 45.127 ;
      RECT 52.037 45.025 54.607 45.081 ;
      RECT 52.083 44.979 54.653 45.035 ;
      RECT 52.129 44.933 54.699 44.989 ;
      RECT 52.175 44.887 54.745 44.943 ;
      RECT 52.221 44.841 54.791 44.897 ;
      RECT 52.267 44.795 54.837 44.851 ;
      RECT 52.313 44.749 54.883 44.805 ;
      RECT 52.359 44.703 54.929 44.759 ;
      RECT 52.405 44.657 54.975 44.713 ;
      RECT 52.451 44.611 55.021 44.667 ;
      RECT 52.497 44.565 55.067 44.621 ;
      RECT 52.543 44.519 55.113 44.575 ;
      RECT 52.589 44.473 55.159 44.529 ;
      RECT 52.635 44.427 55.205 44.483 ;
      RECT 52.681 44.381 55.251 44.437 ;
      RECT 52.727 44.335 55.297 44.391 ;
      RECT 52.773 44.289 55.343 44.345 ;
      RECT 52.819 44.243 55.389 44.299 ;
      RECT 52.865 44.197 55.435 44.253 ;
      RECT 52.911 44.151 55.481 44.207 ;
      RECT 52.957 44.105 55.527 44.161 ;
      RECT 53.003 44.059 55.573 44.115 ;
      RECT 53.049 44.013 55.619 44.069 ;
      RECT 53.095 43.967 55.665 44.023 ;
      RECT 53.141 43.921 55.711 43.977 ;
      RECT 53.187 43.875 55.757 43.931 ;
      RECT 53.233 43.829 55.803 43.885 ;
      RECT 53.279 43.783 55.849 43.839 ;
      RECT 53.325 43.737 55.895 43.793 ;
      RECT 53.371 43.691 55.941 43.747 ;
      RECT 53.417 43.645 55.987 43.701 ;
      RECT 53.463 43.599 56.033 43.655 ;
      RECT 53.509 43.553 56.079 43.609 ;
      RECT 53.555 43.507 56.125 43.563 ;
      RECT 53.601 43.461 56.171 43.517 ;
      RECT 53.647 43.415 56.217 43.471 ;
      RECT 53.693 43.369 56.263 43.425 ;
      RECT 53.739 43.323 56.309 43.379 ;
      RECT 53.785 43.277 56.355 43.333 ;
      RECT 53.831 43.231 56.401 43.287 ;
      RECT 53.877 43.185 56.447 43.241 ;
      RECT 53.923 43.139 56.493 43.195 ;
      RECT 53.969 43.093 56.539 43.149 ;
      RECT 54.015 43.047 56.585 43.103 ;
      RECT 54.061 43.001 56.631 43.057 ;
      RECT 54.107 42.955 56.677 43.011 ;
      RECT 54.153 42.909 56.723 42.965 ;
      RECT 54.199 42.863 56.769 42.919 ;
      RECT 54.245 42.817 56.815 42.873 ;
      RECT 54.291 42.771 56.861 42.827 ;
      RECT 54.337 42.725 56.907 42.781 ;
      RECT 54.383 42.679 56.953 42.735 ;
      RECT 54.429 42.633 56.999 42.689 ;
      RECT 54.475 42.587 57.045 42.643 ;
      RECT 54.521 42.541 57.091 42.597 ;
      RECT 54.567 42.495 57.137 42.551 ;
      RECT 54.613 42.449 57.183 42.505 ;
      RECT 54.659 42.403 57.229 42.459 ;
      RECT 54.705 42.357 57.275 42.413 ;
      RECT 54.751 42.311 57.321 42.367 ;
      RECT 54.797 42.265 57.367 42.321 ;
      RECT 54.843 42.219 57.413 42.275 ;
      RECT 54.889 42.173 57.459 42.229 ;
      RECT 54.935 42.127 57.505 42.183 ;
      RECT 54.981 42.081 57.551 42.137 ;
      RECT 55.027 42.035 57.597 42.091 ;
      RECT 55.073 41.989 57.643 42.045 ;
      RECT 55.119 41.943 57.689 41.999 ;
      RECT 55.165 41.897 57.735 41.953 ;
      RECT 55.211 41.851 57.781 41.907 ;
      RECT 55.257 41.805 57.827 41.861 ;
      RECT 55.303 41.759 57.873 41.815 ;
      RECT 55.349 41.713 57.919 41.769 ;
      RECT 55.395 41.667 57.965 41.723 ;
      RECT 55.441 41.621 58.011 41.677 ;
      RECT 55.487 41.575 58.057 41.631 ;
      RECT 55.533 41.529 58.103 41.585 ;
      RECT 55.579 41.483 58.149 41.539 ;
      RECT 55.625 41.437 58.195 41.493 ;
      RECT 55.671 41.391 58.241 41.447 ;
      RECT 55.717 41.345 58.287 41.401 ;
      RECT 55.763 41.299 58.333 41.355 ;
      RECT 55.809 41.253 58.379 41.309 ;
      RECT 55.855 41.207 58.425 41.263 ;
      RECT 55.901 41.161 58.471 41.217 ;
      RECT 55.947 41.115 58.517 41.171 ;
      RECT 55.993 41.069 58.563 41.125 ;
      RECT 56.039 41.023 58.609 41.079 ;
      RECT 56.085 40.977 58.655 41.033 ;
      RECT 56.131 40.931 58.701 40.987 ;
      RECT 56.177 40.885 58.747 40.941 ;
      RECT 56.223 40.839 58.793 40.895 ;
      RECT 56.269 40.793 58.839 40.849 ;
      RECT 56.315 40.747 58.885 40.803 ;
      RECT 56.361 40.701 58.931 40.757 ;
      RECT 56.407 40.655 58.977 40.711 ;
      RECT 56.453 40.609 59.023 40.665 ;
      RECT 56.499 40.563 59.069 40.619 ;
      RECT 56.545 40.517 59.115 40.573 ;
      RECT 56.591 40.471 59.161 40.527 ;
      RECT 56.637 40.425 59.207 40.481 ;
      RECT 56.683 40.379 59.253 40.435 ;
      RECT 56.729 40.333 59.299 40.389 ;
      RECT 56.775 40.287 59.345 40.343 ;
      RECT 56.821 40.241 59.391 40.297 ;
      RECT 56.867 40.195 59.437 40.251 ;
      RECT 56.913 40.149 59.483 40.205 ;
      RECT 56.959 40.103 59.529 40.159 ;
      RECT 57.005 40.057 59.575 40.113 ;
      RECT 57.051 40.011 59.621 40.067 ;
      RECT 57.097 39.965 59.667 40.021 ;
      RECT 57.143 39.919 59.713 39.975 ;
      RECT 57.189 39.873 59.759 39.929 ;
      RECT 57.235 39.827 59.805 39.883 ;
      RECT 57.281 39.781 59.851 39.837 ;
      RECT 57.327 39.735 59.897 39.791 ;
      RECT 57.373 39.689 59.943 39.745 ;
      RECT 57.419 39.643 59.989 39.699 ;
      RECT 57.465 39.597 60.035 39.653 ;
      RECT 57.511 39.551 60.081 39.607 ;
      RECT 57.557 39.505 60.127 39.561 ;
      RECT 57.603 39.459 60.173 39.515 ;
      RECT 57.649 39.413 60.219 39.469 ;
      RECT 57.695 39.367 60.265 39.423 ;
      RECT 57.741 39.321 60.311 39.377 ;
      RECT 57.787 39.275 60.357 39.331 ;
      RECT 57.833 39.229 60.403 39.285 ;
      RECT 57.879 39.183 60.449 39.239 ;
      RECT 57.925 39.137 60.495 39.193 ;
      RECT 57.971 39.091 60.541 39.147 ;
      RECT 58.017 39.045 60.587 39.101 ;
      RECT 58.063 38.999 60.633 39.055 ;
      RECT 58.109 38.953 60.679 39.009 ;
      RECT 58.155 38.907 60.725 38.963 ;
      RECT 58.201 38.861 60.771 38.917 ;
      RECT 58.247 38.815 60.817 38.871 ;
      RECT 58.293 38.769 60.863 38.825 ;
      RECT 58.339 38.723 60.909 38.779 ;
      RECT 58.385 38.677 60.955 38.733 ;
      RECT 58.431 38.631 61.001 38.687 ;
      RECT 58.477 38.585 61.047 38.641 ;
      RECT 58.523 38.539 61.093 38.595 ;
      RECT 58.569 38.493 61.139 38.549 ;
      RECT 58.615 38.447 61.185 38.503 ;
      RECT 58.661 38.401 61.231 38.457 ;
      RECT 58.707 38.355 61.277 38.411 ;
      RECT 58.753 38.309 61.323 38.365 ;
      RECT 58.799 38.263 61.369 38.319 ;
      RECT 58.845 38.217 61.415 38.273 ;
      RECT 58.891 38.171 61.461 38.227 ;
      RECT 58.937 38.125 61.507 38.181 ;
      RECT 58.983 38.079 61.553 38.135 ;
      RECT 59.029 38.033 61.599 38.089 ;
      RECT 59.075 37.987 61.645 38.043 ;
      RECT 59.121 37.941 61.691 37.997 ;
      RECT 59.167 37.895 61.737 37.951 ;
      RECT 59.213 37.849 61.783 37.905 ;
      RECT 59.259 37.803 61.829 37.859 ;
      RECT 59.305 37.757 61.875 37.813 ;
      RECT 59.351 37.711 61.921 37.767 ;
      RECT 59.397 37.665 61.967 37.721 ;
      RECT 59.443 37.619 62.013 37.675 ;
      RECT 59.489 37.573 62.059 37.629 ;
      RECT 59.535 37.527 62.105 37.583 ;
      RECT 59.581 37.481 62.151 37.537 ;
      RECT 59.627 37.435 62.197 37.491 ;
      RECT 59.673 37.389 62.243 37.445 ;
      RECT 59.719 37.343 62.289 37.399 ;
      RECT 59.765 37.297 62.335 37.353 ;
      RECT 59.811 37.251 62.381 37.307 ;
      RECT 59.857 37.205 62.427 37.261 ;
      RECT 59.903 37.159 62.473 37.215 ;
      RECT 59.949 37.113 62.519 37.169 ;
      RECT 59.995 37.067 62.565 37.123 ;
      RECT 60.041 37.021 62.611 37.077 ;
      RECT 60.087 36.975 62.657 37.031 ;
      RECT 60.133 36.929 62.703 36.985 ;
      RECT 60.179 36.883 62.749 36.939 ;
      RECT 60.225 36.837 62.795 36.893 ;
      RECT 60.271 36.791 62.841 36.847 ;
      RECT 60.317 36.745 62.887 36.801 ;
      RECT 60.363 36.699 62.933 36.755 ;
      RECT 60.409 36.653 62.979 36.709 ;
      RECT 62.939 34.146 62.979 36.709 ;
      RECT 60.455 36.607 63.025 36.663 ;
      RECT 62.94 34.122 63.025 36.663 ;
      RECT 60.501 36.561 63.071 36.617 ;
      RECT 62.986 34.076 63.071 36.617 ;
      RECT 60.547 36.515 63.117 36.571 ;
      RECT 63.032 34.03 63.117 36.571 ;
      RECT 60.593 36.469 63.163 36.525 ;
      RECT 63.078 33.984 63.163 36.525 ;
      RECT 60.639 36.423 63.209 36.479 ;
      RECT 63.124 33.938 63.209 36.479 ;
      RECT 60.685 36.377 63.255 36.433 ;
      RECT 63.17 33.892 63.255 36.433 ;
      RECT 60.731 36.331 63.301 36.387 ;
      RECT 63.216 33.846 63.301 36.387 ;
      RECT 60.777 36.285 63.347 36.341 ;
      RECT 63.262 33.8 63.347 36.341 ;
      RECT 60.823 36.239 63.393 36.295 ;
      RECT 63.308 33.754 63.393 36.295 ;
      RECT 60.869 36.193 63.439 36.249 ;
      RECT 63.354 33.708 63.439 36.249 ;
      RECT 60.915 36.147 63.485 36.203 ;
      RECT 63.4 33.662 63.485 36.203 ;
      RECT 60.961 36.101 63.531 36.157 ;
      RECT 63.446 33.616 63.531 36.157 ;
      RECT 61.007 36.055 63.577 36.111 ;
      RECT 63.492 33.57 63.577 36.111 ;
      RECT 61.053 36.009 63.623 36.065 ;
      RECT 63.538 33.524 63.623 36.065 ;
      RECT 61.099 35.963 63.669 36.019 ;
      RECT 63.584 33.478 63.669 36.019 ;
      RECT 61.145 35.917 63.715 35.973 ;
      RECT 63.63 33.432 63.715 35.973 ;
      RECT 61.191 35.871 63.761 35.927 ;
      RECT 63.676 33.386 63.761 35.927 ;
      RECT 61.237 35.825 63.807 35.881 ;
      RECT 63.722 33.34 63.807 35.881 ;
      RECT 61.283 35.779 63.853 35.835 ;
      RECT 63.768 33.294 63.853 35.835 ;
      RECT 61.329 35.733 63.899 35.789 ;
      RECT 63.814 33.248 63.899 35.789 ;
      RECT 61.375 35.687 63.945 35.743 ;
      RECT 63.86 33.202 63.945 35.743 ;
      RECT 61.421 35.641 63.991 35.697 ;
      RECT 63.906 33.156 63.991 35.697 ;
      RECT 61.467 35.595 64.037 35.651 ;
      RECT 63.952 33.11 64.037 35.651 ;
      RECT 61.513 35.549 64.083 35.605 ;
      RECT 63.998 33.064 64.083 35.605 ;
      RECT 61.559 35.503 64.129 35.559 ;
      RECT 64.044 33.018 64.129 35.559 ;
      RECT 61.605 35.457 64.175 35.513 ;
      RECT 64.09 32.972 64.175 35.513 ;
      RECT 61.651 35.411 64.221 35.467 ;
      RECT 64.136 32.926 64.221 35.467 ;
      RECT 61.697 35.365 64.267 35.421 ;
      RECT 64.182 32.88 64.267 35.421 ;
      RECT 61.743 35.319 64.313 35.375 ;
      RECT 64.228 32.834 64.313 35.375 ;
      RECT 61.789 35.273 64.359 35.329 ;
      RECT 64.274 32.788 64.359 35.329 ;
      RECT 61.835 35.227 64.405 35.283 ;
      RECT 64.32 32.742 64.405 35.283 ;
      RECT 61.881 35.181 64.451 35.237 ;
      RECT 64.366 32.696 64.451 35.237 ;
      RECT 61.927 35.135 64.497 35.191 ;
      RECT 64.412 32.65 64.497 35.191 ;
      RECT 61.973 35.089 64.543 35.145 ;
      RECT 64.458 32.604 64.543 35.145 ;
      RECT 62.019 35.043 64.589 35.099 ;
      RECT 64.504 32.558 64.589 35.099 ;
      RECT 62.065 34.997 64.635 35.053 ;
      RECT 64.55 32.512 64.635 35.053 ;
      RECT 62.111 34.951 64.681 35.007 ;
      RECT 64.596 32.466 64.681 35.007 ;
      RECT 62.157 34.905 64.727 34.961 ;
      RECT 64.642 32.42 64.727 34.961 ;
      RECT 62.203 34.859 64.773 34.915 ;
      RECT 64.688 32.374 64.773 34.915 ;
      RECT 62.249 34.813 64.819 34.869 ;
      RECT 64.734 32.328 64.819 34.869 ;
      RECT 62.295 34.767 64.865 34.823 ;
      RECT 64.78 32.282 64.865 34.823 ;
      RECT 62.341 34.721 64.911 34.777 ;
      RECT 64.826 32.236 64.911 34.777 ;
      RECT 62.387 34.675 64.957 34.731 ;
      RECT 64.872 32.19 64.957 34.731 ;
      RECT 62.433 34.629 65.003 34.685 ;
      RECT 64.918 32.144 65.003 34.685 ;
      RECT 62.479 34.583 65.049 34.639 ;
      RECT 64.964 32.098 65.049 34.639 ;
      RECT 62.525 34.537 65.095 34.593 ;
      RECT 65.01 32.052 65.095 34.593 ;
      RECT 62.571 34.491 65.141 34.547 ;
      RECT 65.056 32.006 65.141 34.547 ;
      RECT 62.617 34.445 65.187 34.501 ;
      RECT 65.102 31.96 65.187 34.501 ;
      RECT 62.663 34.399 65.233 34.455 ;
      RECT 65.148 31.914 65.233 34.455 ;
      RECT 62.709 34.353 65.279 34.409 ;
      RECT 65.194 31.868 65.279 34.409 ;
      RECT 62.755 34.307 65.325 34.363 ;
      RECT 65.24 31.822 65.325 34.363 ;
      RECT 62.801 34.261 65.371 34.317 ;
      RECT 65.286 31.776 65.371 34.317 ;
      RECT 62.847 34.215 65.417 34.271 ;
      RECT 65.332 31.73 65.417 34.271 ;
      RECT 62.893 34.169 65.463 34.225 ;
      RECT 65.378 31.684 65.463 34.225 ;
      RECT 65.424 31.638 65.509 34.179 ;
      RECT 65.47 31.592 65.555 34.133 ;
      RECT 65.516 31.546 65.601 34.087 ;
      RECT 65.562 31.5 65.647 34.041 ;
      RECT 65.608 31.454 65.693 33.995 ;
      RECT 65.654 31.408 65.739 33.949 ;
      RECT 65.7 31.362 65.785 33.903 ;
      RECT 65.746 31.316 65.831 33.857 ;
      RECT 65.792 31.27 65.877 33.811 ;
      RECT 65.838 31.224 65.923 33.765 ;
      RECT 65.884 31.178 65.969 33.719 ;
      RECT 65.93 31.132 66.015 33.673 ;
      RECT 65.976 31.086 66.061 33.627 ;
      RECT 66.022 31.04 66.107 33.581 ;
      RECT 66.068 30.994 66.153 33.535 ;
      RECT 66.114 30.948 66.199 33.489 ;
      RECT 66.16 30.902 66.245 33.443 ;
      RECT 66.206 30.856 66.291 33.397 ;
      RECT 66.252 30.81 66.337 33.351 ;
      RECT 66.298 30.764 66.383 33.305 ;
      RECT 66.344 30.718 66.429 33.259 ;
      RECT 66.39 30.672 66.475 33.213 ;
      RECT 66.436 30.626 66.521 33.167 ;
      RECT 66.482 30.58 66.567 33.121 ;
      RECT 66.528 30.534 66.613 33.075 ;
      RECT 66.574 30.488 66.659 33.029 ;
      RECT 66.62 30.442 66.705 32.983 ;
      RECT 66.666 30.396 66.751 32.937 ;
      RECT 66.712 30.35 66.797 32.891 ;
      RECT 66.758 30.304 66.843 32.845 ;
      RECT 66.804 30.258 66.889 32.799 ;
      RECT 66.85 30.212 66.935 32.753 ;
      RECT 66.896 30.166 66.981 32.707 ;
      RECT 66.942 30.12 67.027 32.661 ;
      RECT 66.988 30.074 67.073 32.615 ;
      RECT 67.034 30.028 67.119 32.569 ;
      RECT 67.08 29.982 67.165 32.523 ;
      RECT 67.126 29.936 67.211 32.477 ;
      RECT 67.172 29.89 67.257 32.431 ;
      RECT 67.218 29.844 67.303 32.385 ;
      RECT 67.264 29.798 67.349 32.339 ;
      RECT 67.31 29.752 67.395 32.293 ;
      RECT 67.356 29.706 67.441 32.247 ;
      RECT 67.402 29.66 67.487 32.201 ;
      RECT 67.448 29.614 67.533 32.155 ;
      RECT 67.494 29.568 67.579 32.109 ;
      RECT 67.54 29.522 67.625 32.063 ;
      RECT 67.586 29.476 67.671 32.017 ;
      RECT 67.632 29.43 67.717 31.971 ;
      RECT 67.678 29.384 67.763 31.925 ;
      RECT 67.724 29.338 67.809 31.879 ;
      RECT 67.77 29.292 67.855 31.833 ;
      RECT 67.816 29.246 67.901 31.787 ;
      RECT 67.862 29.199 67.947 31.741 ;
      RECT 67.908 29.175 67.993 31.695 ;
      RECT 67.908 29.175 68.039 31.649 ;
      RECT 67.908 29.175 68.085 31.603 ;
      RECT 67.908 29.175 68.131 31.557 ;
      RECT 67.908 29.175 68.177 31.511 ;
      RECT 67.908 29.175 68.223 31.465 ;
      RECT 67.908 29.175 68.269 31.419 ;
      RECT 67.908 29.175 68.315 31.373 ;
      RECT 67.908 29.175 68.361 31.327 ;
      RECT 67.908 29.175 68.407 31.281 ;
      RECT 67.908 29.175 68.453 31.235 ;
      RECT 67.908 29.175 68.499 31.189 ;
      RECT 67.908 29.175 68.545 31.143 ;
      RECT 67.908 29.175 68.591 31.097 ;
      RECT 67.908 29.175 68.637 31.051 ;
      RECT 67.908 29.175 68.683 31.005 ;
      RECT 67.908 29.175 68.729 30.959 ;
      RECT 67.908 29.175 68.775 30.913 ;
      RECT 67.908 29.175 68.821 30.867 ;
      RECT 67.908 29.175 68.867 30.821 ;
      RECT 67.908 29.175 68.913 30.775 ;
      RECT 67.908 29.175 68.959 30.729 ;
      RECT 67.908 29.175 69.005 30.683 ;
      RECT 67.908 29.175 69.051 30.637 ;
      RECT 67.908 29.175 69.097 30.591 ;
      RECT 67.908 29.175 69.143 30.545 ;
      RECT 67.908 29.175 69.189 30.499 ;
      RECT 67.908 29.175 69.235 30.453 ;
      RECT 67.908 29.175 69.281 30.407 ;
      RECT 67.908 29.175 69.327 30.361 ;
      RECT 66.758 30.304 69.34 30.331 ;
      RECT 67.908 29.175 110 30.325 ;
      RECT 42.675 74.637 43.825 110 ;
      RECT 42.675 74.637 43.871 76.067 ;
      RECT 42.675 74.637 43.917 76.021 ;
      RECT 42.675 74.637 43.963 75.975 ;
      RECT 42.675 74.637 44.009 75.929 ;
      RECT 42.675 74.637 44.055 75.883 ;
      RECT 42.675 74.637 44.101 75.837 ;
      RECT 42.675 74.637 44.147 75.791 ;
      RECT 42.675 74.637 44.193 75.745 ;
      RECT 42.675 74.637 44.239 75.699 ;
      RECT 42.675 74.637 44.285 75.653 ;
      RECT 42.675 74.637 44.331 75.607 ;
      RECT 42.675 74.637 44.377 75.561 ;
      RECT 42.675 74.637 44.423 75.515 ;
      RECT 42.675 74.637 44.469 75.469 ;
      RECT 42.675 74.637 44.515 75.423 ;
      RECT 42.675 74.637 44.561 75.377 ;
      RECT 42.675 74.637 44.607 75.331 ;
      RECT 42.675 74.637 44.653 75.285 ;
      RECT 42.675 74.637 44.699 75.239 ;
      RECT 42.675 74.637 44.745 75.193 ;
      RECT 42.675 74.637 44.791 75.147 ;
      RECT 42.675 74.637 44.837 75.101 ;
      RECT 42.675 74.637 44.883 75.055 ;
      RECT 42.675 74.637 44.929 75.009 ;
      RECT 42.675 74.637 44.975 74.963 ;
      RECT 42.675 74.637 45.021 74.917 ;
      RECT 42.675 74.637 45.067 74.871 ;
      RECT 42.675 74.637 45.113 74.825 ;
      RECT 42.675 74.637 45.159 74.779 ;
      RECT 42.675 74.637 45.205 74.733 ;
      RECT 42.675 74.637 45.251 74.687 ;
      RECT 42.721 74.591 45.297 74.641 ;
      RECT 42.767 74.545 45.343 74.595 ;
      RECT 42.813 74.499 45.389 74.549 ;
      RECT 42.859 74.453 45.435 74.503 ;
      RECT 42.905 74.407 45.481 74.457 ;
      RECT 42.951 74.361 45.527 74.411 ;
      RECT 42.997 74.315 45.573 74.365 ;
      RECT 43.043 74.269 45.619 74.319 ;
      RECT 43.089 74.223 45.665 74.273 ;
      RECT 43.135 74.177 45.711 74.227 ;
      RECT 43.181 74.131 45.757 74.181 ;
      RECT 43.227 74.085 45.803 74.135 ;
      RECT 43.273 74.039 45.849 74.089 ;
      RECT 43.319 73.993 45.895 74.043 ;
      RECT 43.365 73.947 45.941 73.997 ;
      RECT 43.411 73.901 45.987 73.951 ;
      RECT 43.457 73.855 46.033 73.905 ;
      RECT 43.503 73.809 46.079 73.859 ;
      RECT 43.549 73.763 46.125 73.813 ;
      RECT 43.595 73.717 46.171 73.767 ;
      RECT 43.641 73.671 46.217 73.721 ;
      RECT 43.687 73.625 46.263 73.675 ;
      RECT 43.733 73.579 46.309 73.629 ;
      RECT 43.779 73.533 46.355 73.583 ;
      RECT 43.825 73.487 46.401 73.537 ;
      RECT 43.871 73.441 46.447 73.491 ;
      RECT 43.917 73.395 46.493 73.445 ;
      RECT 43.963 73.349 46.539 73.399 ;
      RECT 44.009 73.303 46.585 73.353 ;
      RECT 44.055 73.257 46.631 73.307 ;
      RECT 44.101 73.211 46.677 73.261 ;
      RECT 44.147 73.165 46.723 73.215 ;
      RECT 44.193 73.119 46.769 73.169 ;
      RECT 44.239 73.073 46.815 73.123 ;
      RECT 44.285 73.027 46.861 73.077 ;
      RECT 44.331 72.981 46.907 73.031 ;
      RECT 44.377 72.935 46.953 72.985 ;
      RECT 44.423 72.889 46.999 72.939 ;
      RECT 44.469 72.843 47.045 72.893 ;
      RECT 44.515 72.797 47.091 72.847 ;
      RECT 44.561 72.751 47.137 72.801 ;
      RECT 44.607 72.705 47.183 72.755 ;
      RECT 44.653 72.659 47.229 72.709 ;
      RECT 44.699 72.613 47.275 72.663 ;
      RECT 44.745 72.567 47.321 72.617 ;
      RECT 44.791 72.521 47.367 72.571 ;
      RECT 44.837 72.475 47.413 72.525 ;
      RECT 44.883 72.429 47.459 72.479 ;
      RECT 44.929 72.383 47.505 72.433 ;
      RECT 44.975 72.337 47.551 72.387 ;
      RECT 45.021 72.291 47.597 72.341 ;
      RECT 45.067 72.245 47.643 72.295 ;
      RECT 45.113 72.199 47.689 72.249 ;
      RECT 45.159 72.153 47.735 72.203 ;
      RECT 45.205 72.107 47.781 72.157 ;
      RECT 45.251 72.061 47.827 72.111 ;
      RECT 45.297 72.015 47.873 72.065 ;
      RECT 45.343 71.969 47.919 72.019 ;
      RECT 45.389 71.923 47.965 71.973 ;
      RECT 45.435 71.877 48.011 71.927 ;
      RECT 45.481 71.831 48.057 71.881 ;
      RECT 45.527 71.785 48.103 71.835 ;
      RECT 45.573 71.739 48.149 71.789 ;
      RECT 45.619 71.693 48.195 71.743 ;
      RECT 45.665 71.647 48.241 71.697 ;
      RECT 45.711 71.601 48.287 71.651 ;
      RECT 45.757 71.555 48.333 71.605 ;
      RECT 45.803 71.509 48.379 71.559 ;
      RECT 45.849 71.463 48.425 71.513 ;
      RECT 45.895 71.417 48.471 71.467 ;
      RECT 45.941 71.371 48.517 71.421 ;
      RECT 45.987 71.325 48.563 71.375 ;
      RECT 46.033 71.279 48.609 71.329 ;
      RECT 46.079 71.233 48.655 71.283 ;
      RECT 46.125 71.187 48.701 71.237 ;
      RECT 46.171 71.141 48.747 71.191 ;
      RECT 46.217 71.095 48.793 71.145 ;
      RECT 46.263 71.049 48.839 71.099 ;
      RECT 46.309 71.003 48.885 71.053 ;
      RECT 46.355 70.957 48.931 71.007 ;
      RECT 46.401 70.911 48.977 70.961 ;
      RECT 46.447 70.865 49.023 70.915 ;
      RECT 46.493 70.819 49.069 70.869 ;
      RECT 46.539 70.773 49.115 70.823 ;
      RECT 46.585 70.727 49.161 70.777 ;
      RECT 46.631 70.681 49.207 70.731 ;
      RECT 46.677 70.635 49.253 70.685 ;
      RECT 46.723 70.589 49.299 70.639 ;
      RECT 46.769 70.543 49.345 70.593 ;
      RECT 46.815 70.497 49.391 70.547 ;
      RECT 46.861 70.451 49.437 70.501 ;
      RECT 46.907 70.405 49.483 70.455 ;
      RECT 46.953 70.359 49.529 70.409 ;
      RECT 46.999 70.313 49.575 70.363 ;
      RECT 47.045 70.267 49.621 70.317 ;
      RECT 47.091 70.221 49.667 70.271 ;
      RECT 47.137 70.175 49.713 70.225 ;
      RECT 47.183 70.129 49.759 70.179 ;
      RECT 47.229 70.083 49.805 70.133 ;
      RECT 47.275 70.037 49.851 70.087 ;
      RECT 47.321 69.991 49.897 70.041 ;
      RECT 47.367 69.945 49.943 69.995 ;
      RECT 47.413 69.899 49.989 69.949 ;
      RECT 47.459 69.853 50.035 69.903 ;
      RECT 47.505 69.807 50.081 69.857 ;
      RECT 47.551 69.761 50.127 69.811 ;
      RECT 47.597 69.715 50.173 69.765 ;
      RECT 47.643 69.669 50.219 69.719 ;
      RECT 47.689 69.623 50.265 69.673 ;
      RECT 47.735 69.577 50.311 69.627 ;
      RECT 47.781 69.531 50.357 69.581 ;
      RECT 47.827 69.485 50.403 69.535 ;
      RECT 47.873 69.439 50.449 69.489 ;
      RECT 47.919 69.393 50.495 69.443 ;
      RECT 47.965 69.347 50.541 69.397 ;
      RECT 48.011 69.301 50.587 69.351 ;
      RECT 48.057 69.255 50.633 69.305 ;
      RECT 48.103 69.209 50.679 69.259 ;
      RECT 48.149 69.163 50.725 69.213 ;
      RECT 48.195 69.117 50.771 69.167 ;
      RECT 48.241 69.071 50.817 69.121 ;
      RECT 48.287 69.025 50.863 69.075 ;
      RECT 48.333 68.979 50.909 69.029 ;
      RECT 48.379 68.933 50.955 68.983 ;
      RECT 48.425 68.887 51.001 68.937 ;
      RECT 48.471 68.841 51.047 68.891 ;
      RECT 48.517 68.795 51.093 68.845 ;
      RECT 48.563 68.749 51.139 68.799 ;
      RECT 48.609 68.703 51.185 68.753 ;
      RECT 48.655 68.657 51.231 68.707 ;
      RECT 48.701 68.611 51.277 68.661 ;
      RECT 48.747 68.565 51.323 68.615 ;
      RECT 48.793 68.519 51.369 68.569 ;
      RECT 48.839 68.473 51.415 68.523 ;
      RECT 48.885 68.427 51.461 68.477 ;
      RECT 48.931 68.381 51.507 68.431 ;
      RECT 48.977 68.335 51.553 68.385 ;
      RECT 49.023 68.289 51.599 68.339 ;
      RECT 49.069 68.243 51.645 68.293 ;
      RECT 49.115 68.197 51.691 68.247 ;
      RECT 49.161 68.151 51.737 68.201 ;
      RECT 49.207 68.105 51.783 68.155 ;
      RECT 49.253 68.059 51.829 68.109 ;
      RECT 49.299 68.013 51.875 68.063 ;
      RECT 49.345 67.967 51.921 68.017 ;
      RECT 49.391 67.921 51.967 67.971 ;
      RECT 49.437 67.875 52.013 67.925 ;
      RECT 49.483 67.829 52.059 67.879 ;
      RECT 49.529 67.783 52.105 67.833 ;
      RECT 49.575 67.737 52.151 67.787 ;
      RECT 49.621 67.691 52.197 67.741 ;
      RECT 49.667 67.645 52.243 67.695 ;
      RECT 49.713 67.599 52.289 67.649 ;
      RECT 49.759 67.553 52.335 67.603 ;
      RECT 49.805 67.507 52.381 67.557 ;
      RECT 49.851 67.461 52.427 67.511 ;
      RECT 49.897 67.415 52.473 67.465 ;
      RECT 49.943 67.369 52.519 67.419 ;
      RECT 49.989 67.323 52.565 67.373 ;
      RECT 50.035 67.277 52.611 67.327 ;
      RECT 50.081 67.231 52.657 67.281 ;
      RECT 50.127 67.185 52.703 67.235 ;
      RECT 50.173 67.139 52.749 67.189 ;
      RECT 50.219 67.093 52.795 67.143 ;
      RECT 50.265 67.047 52.841 67.097 ;
      RECT 50.311 67.001 52.887 67.051 ;
      RECT 50.357 66.955 52.933 67.005 ;
      RECT 50.403 66.909 52.979 66.959 ;
      RECT 50.449 66.863 53.025 66.913 ;
      RECT 50.495 66.817 53.071 66.867 ;
      RECT 50.541 66.771 53.117 66.821 ;
      RECT 50.587 66.725 53.163 66.775 ;
      RECT 50.633 66.679 53.209 66.729 ;
      RECT 50.679 66.633 53.255 66.683 ;
      RECT 50.725 66.587 53.301 66.637 ;
      RECT 50.771 66.541 53.347 66.591 ;
      RECT 50.817 66.495 53.393 66.545 ;
      RECT 50.863 66.449 53.439 66.499 ;
      RECT 50.909 66.403 53.485 66.453 ;
      RECT 50.955 66.357 53.531 66.407 ;
      RECT 51.001 66.311 53.577 66.361 ;
      RECT 51.047 66.265 53.623 66.315 ;
      RECT 51.093 66.219 53.669 66.269 ;
      RECT 51.139 66.173 53.715 66.223 ;
      RECT 51.185 66.127 53.761 66.177 ;
      RECT 51.231 66.081 53.807 66.131 ;
      RECT 51.277 66.035 53.853 66.085 ;
      RECT 51.323 65.989 53.899 66.039 ;
      RECT 51.369 65.943 53.945 65.993 ;
      RECT 51.415 65.897 53.991 65.947 ;
      RECT 51.461 65.851 54.037 65.901 ;
      RECT 51.507 65.805 54.083 65.855 ;
      RECT 51.553 65.759 54.129 65.809 ;
      RECT 51.599 65.713 54.175 65.763 ;
      RECT 51.645 65.667 54.221 65.717 ;
      RECT 51.691 65.621 54.267 65.671 ;
      RECT 51.737 65.575 54.313 65.625 ;
      RECT 51.783 65.529 54.359 65.579 ;
      RECT 51.829 65.483 54.405 65.533 ;
      RECT 51.875 65.437 54.451 65.487 ;
      RECT 51.921 65.391 54.497 65.441 ;
      RECT 51.967 65.345 54.543 65.395 ;
      RECT 52.013 65.299 54.589 65.349 ;
      RECT 52.059 65.253 54.635 65.303 ;
      RECT 52.105 65.207 54.681 65.257 ;
      RECT 52.151 65.161 54.727 65.211 ;
      RECT 52.197 65.115 54.773 65.165 ;
      RECT 52.243 65.069 54.819 65.119 ;
      RECT 52.289 65.023 54.865 65.073 ;
      RECT 52.335 64.977 54.911 65.027 ;
      RECT 52.381 64.931 54.957 64.981 ;
      RECT 52.427 64.885 55.003 64.935 ;
      RECT 52.473 64.839 55.049 64.889 ;
      RECT 52.519 64.793 55.095 64.843 ;
      RECT 52.565 64.747 55.141 64.797 ;
      RECT 52.611 64.701 55.187 64.751 ;
      RECT 52.657 64.655 55.233 64.705 ;
      RECT 52.703 64.609 55.279 64.659 ;
      RECT 52.749 64.563 55.325 64.613 ;
      RECT 52.795 64.517 55.371 64.567 ;
      RECT 52.841 64.471 55.417 64.521 ;
      RECT 52.887 64.425 55.463 64.475 ;
      RECT 52.933 64.379 55.509 64.429 ;
      RECT 52.979 64.333 55.555 64.383 ;
      RECT 53.025 64.287 55.601 64.337 ;
      RECT 53.071 64.241 55.647 64.291 ;
      RECT 53.117 64.195 55.693 64.245 ;
      RECT 53.163 64.149 55.739 64.199 ;
      RECT 53.209 64.103 55.785 64.153 ;
      RECT 53.255 64.057 55.825 64.11 ;
      RECT 53.301 64.011 55.871 64.067 ;
      RECT 53.347 63.965 55.917 64.021 ;
      RECT 53.393 63.919 55.963 63.975 ;
      RECT 53.439 63.873 56.009 63.929 ;
      RECT 53.485 63.827 56.055 63.883 ;
      RECT 53.531 63.781 56.101 63.837 ;
      RECT 53.577 63.735 56.147 63.791 ;
      RECT 53.623 63.689 56.193 63.745 ;
      RECT 53.669 63.643 56.239 63.699 ;
      RECT 53.715 63.597 56.285 63.653 ;
      RECT 53.761 63.551 56.331 63.607 ;
      RECT 53.807 63.505 56.377 63.561 ;
      RECT 53.853 63.459 56.423 63.515 ;
      RECT 53.899 63.413 56.469 63.469 ;
      RECT 53.945 63.367 56.515 63.423 ;
      RECT 53.991 63.321 56.561 63.377 ;
      RECT 54.037 63.275 56.607 63.331 ;
      RECT 54.083 63.229 56.653 63.285 ;
      RECT 54.129 63.183 56.699 63.239 ;
      RECT 54.175 63.137 56.745 63.193 ;
      RECT 54.221 63.091 56.791 63.147 ;
      RECT 54.267 63.045 56.837 63.101 ;
      RECT 54.313 62.999 56.883 63.055 ;
      RECT 54.359 62.953 56.929 63.009 ;
      RECT 54.405 62.907 56.975 62.963 ;
      RECT 54.451 62.861 57.021 62.917 ;
      RECT 54.497 62.815 57.067 62.871 ;
      RECT 54.543 62.769 57.113 62.825 ;
      RECT 54.589 62.723 57.159 62.779 ;
      RECT 54.635 62.677 57.205 62.733 ;
      RECT 54.681 62.631 57.251 62.687 ;
      RECT 54.727 62.585 57.297 62.641 ;
      RECT 54.773 62.539 57.343 62.595 ;
      RECT 54.819 62.493 57.389 62.549 ;
      RECT 54.865 62.447 57.435 62.503 ;
      RECT 54.911 62.401 57.481 62.457 ;
      RECT 54.957 62.355 57.527 62.411 ;
      RECT 55.003 62.309 57.573 62.365 ;
      RECT 55.049 62.263 57.619 62.319 ;
      RECT 55.095 62.217 57.665 62.273 ;
      RECT 55.141 62.171 57.711 62.227 ;
      RECT 55.187 62.125 57.757 62.181 ;
      RECT 55.233 62.079 57.803 62.135 ;
      RECT 55.279 62.033 57.849 62.089 ;
      RECT 55.325 61.987 57.895 62.043 ;
      RECT 55.371 61.941 57.941 61.997 ;
      RECT 55.417 61.895 57.987 61.951 ;
      RECT 55.463 61.849 58.033 61.905 ;
      RECT 55.509 61.803 58.079 61.859 ;
      RECT 55.555 61.757 58.125 61.813 ;
      RECT 55.601 61.711 58.171 61.767 ;
      RECT 55.647 61.665 58.217 61.721 ;
      RECT 55.693 61.619 58.263 61.675 ;
      RECT 55.739 61.573 58.309 61.629 ;
      RECT 55.785 61.527 58.355 61.583 ;
      RECT 55.831 61.481 58.401 61.537 ;
      RECT 55.877 61.435 58.447 61.491 ;
      RECT 55.923 61.389 58.493 61.445 ;
      RECT 55.969 61.343 58.539 61.399 ;
      RECT 56.015 61.297 58.585 61.353 ;
      RECT 56.061 61.251 58.631 61.307 ;
      RECT 56.107 61.205 58.677 61.261 ;
      RECT 56.153 61.159 58.723 61.215 ;
      RECT 56.199 61.113 58.769 61.169 ;
      RECT 56.245 61.067 58.815 61.123 ;
      RECT 56.291 61.021 58.861 61.077 ;
      RECT 56.337 60.975 58.907 61.031 ;
      RECT 56.383 60.929 58.953 60.985 ;
      RECT 56.429 60.883 58.999 60.939 ;
      RECT 56.475 60.837 59.045 60.893 ;
      RECT 56.521 60.791 59.091 60.847 ;
      RECT 56.567 60.745 59.137 60.801 ;
      RECT 56.613 60.699 59.183 60.755 ;
      RECT 56.659 60.653 59.229 60.709 ;
      RECT 56.705 60.607 59.275 60.663 ;
      RECT 56.751 60.561 59.321 60.617 ;
      RECT 56.797 60.515 59.367 60.571 ;
      RECT 56.843 60.469 59.413 60.525 ;
      RECT 56.889 60.423 59.459 60.479 ;
      RECT 56.935 60.377 59.505 60.433 ;
      RECT 56.981 60.331 59.551 60.387 ;
      RECT 57.027 60.285 59.597 60.341 ;
      RECT 57.073 60.239 59.643 60.295 ;
      RECT 57.119 60.193 59.689 60.249 ;
      RECT 57.165 60.147 59.735 60.203 ;
      RECT 57.211 60.101 59.781 60.157 ;
      RECT 57.257 60.055 59.827 60.111 ;
      RECT 57.303 60.009 59.873 60.065 ;
      RECT 57.349 59.963 59.919 60.019 ;
      RECT 57.395 59.917 59.965 59.973 ;
      RECT 57.441 59.871 60.011 59.927 ;
      RECT 57.487 59.825 60.057 59.881 ;
      RECT 57.533 59.779 60.103 59.835 ;
      RECT 57.579 59.733 60.149 59.789 ;
      RECT 57.625 59.687 60.195 59.743 ;
      RECT 57.671 59.641 60.241 59.697 ;
      RECT 57.717 59.595 60.287 59.651 ;
      RECT 57.763 59.549 60.333 59.605 ;
      RECT 57.809 59.503 60.379 59.559 ;
      RECT 57.855 59.457 60.425 59.513 ;
      RECT 57.901 59.411 60.471 59.467 ;
      RECT 57.947 59.365 60.517 59.421 ;
      RECT 57.993 59.319 60.563 59.375 ;
      RECT 58.039 59.273 60.609 59.329 ;
      RECT 58.085 59.227 60.655 59.283 ;
      RECT 58.131 59.181 60.701 59.237 ;
      RECT 58.177 59.135 60.747 59.191 ;
      RECT 58.223 59.089 60.793 59.145 ;
      RECT 58.269 59.043 60.839 59.099 ;
      RECT 58.315 58.997 60.885 59.053 ;
      RECT 58.361 58.951 60.931 59.007 ;
      RECT 58.407 58.905 60.977 58.961 ;
      RECT 58.453 58.859 61.023 58.915 ;
      RECT 58.499 58.813 61.069 58.869 ;
      RECT 58.545 58.767 61.115 58.823 ;
      RECT 58.591 58.721 61.161 58.777 ;
      RECT 58.637 58.675 61.207 58.731 ;
      RECT 58.683 58.629 61.253 58.685 ;
      RECT 58.729 58.583 61.299 58.639 ;
      RECT 58.775 58.537 61.345 58.593 ;
      RECT 58.821 58.491 61.391 58.547 ;
      RECT 58.867 58.445 61.437 58.501 ;
      RECT 58.913 58.399 61.483 58.455 ;
      RECT 58.959 58.353 61.529 58.409 ;
      RECT 59.005 58.307 61.575 58.363 ;
      RECT 59.051 58.261 61.621 58.317 ;
      RECT 59.097 58.215 61.667 58.271 ;
      RECT 59.143 58.169 61.713 58.225 ;
      RECT 59.189 58.123 61.759 58.179 ;
      RECT 59.235 58.077 61.805 58.133 ;
      RECT 59.281 58.031 61.851 58.087 ;
      RECT 59.327 57.985 61.897 58.041 ;
      RECT 59.373 57.939 61.943 57.995 ;
      RECT 59.419 57.893 61.989 57.949 ;
      RECT 59.465 57.847 62.035 57.903 ;
      RECT 59.511 57.801 62.081 57.857 ;
      RECT 59.557 57.755 62.127 57.811 ;
      RECT 59.603 57.709 62.173 57.765 ;
      RECT 59.649 57.663 62.219 57.719 ;
      RECT 59.695 57.617 62.265 57.673 ;
      RECT 59.741 57.571 62.311 57.627 ;
      RECT 59.787 57.525 62.357 57.581 ;
      RECT 59.833 57.479 62.403 57.535 ;
      RECT 59.879 57.433 62.449 57.489 ;
      RECT 59.925 57.387 62.495 57.443 ;
      RECT 59.971 57.341 62.541 57.397 ;
      RECT 60.017 57.295 62.587 57.351 ;
      RECT 60.063 57.249 62.633 57.305 ;
      RECT 60.109 57.203 62.679 57.259 ;
      RECT 60.155 57.157 62.725 57.213 ;
      RECT 60.201 57.111 62.771 57.167 ;
      RECT 60.247 57.065 62.817 57.121 ;
      RECT 60.293 57.019 62.863 57.075 ;
      RECT 60.339 56.973 62.909 57.029 ;
      RECT 60.385 56.927 62.955 56.983 ;
      RECT 60.431 56.881 63.001 56.937 ;
      RECT 60.477 56.835 63.047 56.891 ;
      RECT 60.523 56.789 63.093 56.845 ;
      RECT 60.569 56.743 63.139 56.799 ;
      RECT 60.615 56.697 63.185 56.753 ;
      RECT 60.661 56.651 63.231 56.707 ;
      RECT 60.707 56.605 63.277 56.661 ;
      RECT 60.753 56.559 63.323 56.615 ;
      RECT 60.799 56.513 63.369 56.569 ;
      RECT 60.845 56.467 63.415 56.523 ;
      RECT 60.891 56.421 63.461 56.477 ;
      RECT 60.937 56.375 63.507 56.431 ;
      RECT 60.983 56.329 63.553 56.385 ;
      RECT 61.029 56.283 63.599 56.339 ;
      RECT 61.075 56.237 63.645 56.293 ;
      RECT 61.121 56.191 63.691 56.247 ;
      RECT 61.167 56.145 63.737 56.201 ;
      RECT 61.213 56.099 63.783 56.155 ;
      RECT 61.259 56.053 63.829 56.109 ;
      RECT 61.305 56.007 63.875 56.063 ;
      RECT 61.351 55.961 63.921 56.017 ;
      RECT 61.397 55.915 63.967 55.971 ;
      RECT 61.443 55.869 64.013 55.925 ;
      RECT 61.489 55.823 64.059 55.879 ;
      RECT 61.535 55.777 64.105 55.833 ;
      RECT 61.581 55.731 64.151 55.787 ;
      RECT 61.627 55.685 64.197 55.741 ;
      RECT 61.673 55.639 64.243 55.695 ;
      RECT 61.719 55.593 64.289 55.649 ;
      RECT 61.765 55.547 64.335 55.603 ;
      RECT 61.811 55.501 64.381 55.557 ;
      RECT 61.857 55.455 64.427 55.511 ;
      RECT 61.903 55.409 64.473 55.465 ;
      RECT 61.949 55.363 64.519 55.419 ;
      RECT 61.995 55.317 64.565 55.373 ;
      RECT 62.041 55.271 64.611 55.327 ;
      RECT 62.087 55.225 64.657 55.281 ;
      RECT 62.133 55.179 64.703 55.235 ;
      RECT 62.179 55.133 64.749 55.189 ;
      RECT 62.225 55.087 64.795 55.143 ;
      RECT 62.271 55.041 64.841 55.097 ;
      RECT 62.317 54.995 64.887 55.051 ;
      RECT 62.363 54.949 64.933 55.005 ;
      RECT 62.409 54.903 64.979 54.959 ;
      RECT 62.455 54.857 65.025 54.913 ;
      RECT 62.501 54.811 65.071 54.867 ;
      RECT 62.547 54.765 65.117 54.821 ;
      RECT 62.593 54.719 65.163 54.775 ;
      RECT 62.639 54.673 65.209 54.729 ;
      RECT 62.685 54.627 65.255 54.683 ;
      RECT 62.731 54.581 65.301 54.637 ;
      RECT 62.777 54.535 65.347 54.591 ;
      RECT 62.823 54.489 65.393 54.545 ;
      RECT 62.869 54.443 65.439 54.499 ;
      RECT 62.915 54.397 65.485 54.453 ;
      RECT 62.961 54.351 65.531 54.407 ;
      RECT 63.007 54.305 65.577 54.361 ;
      RECT 63.053 54.259 65.623 54.315 ;
      RECT 63.099 54.213 65.669 54.269 ;
      RECT 63.145 54.167 65.715 54.223 ;
      RECT 63.191 54.121 65.761 54.177 ;
      RECT 63.237 54.075 65.807 54.131 ;
      RECT 63.283 54.029 65.853 54.085 ;
      RECT 63.329 53.983 65.899 54.039 ;
      RECT 63.375 53.937 65.945 53.993 ;
      RECT 63.421 53.891 65.991 53.947 ;
      RECT 63.467 53.845 66.037 53.901 ;
      RECT 63.513 53.799 66.083 53.855 ;
      RECT 63.559 53.753 66.129 53.809 ;
      RECT 63.605 53.707 66.175 53.763 ;
      RECT 63.651 53.661 66.221 53.717 ;
      RECT 63.697 53.615 66.267 53.671 ;
      RECT 63.743 53.569 66.313 53.625 ;
      RECT 63.789 53.523 66.359 53.579 ;
      RECT 63.835 53.477 66.405 53.533 ;
      RECT 63.881 53.431 66.451 53.487 ;
      RECT 63.927 53.385 66.497 53.441 ;
      RECT 63.973 53.339 66.543 53.395 ;
      RECT 64.019 53.293 66.589 53.349 ;
      RECT 64.065 53.247 66.635 53.303 ;
      RECT 64.111 53.201 66.681 53.257 ;
      RECT 64.157 53.155 66.727 53.211 ;
      RECT 64.203 53.109 66.773 53.165 ;
      RECT 64.249 53.063 66.819 53.119 ;
      RECT 64.295 53.017 66.865 53.073 ;
      RECT 64.341 52.971 66.911 53.027 ;
      RECT 64.387 52.925 66.957 52.981 ;
      RECT 64.433 52.879 67.003 52.935 ;
      RECT 64.479 52.833 67.049 52.889 ;
      RECT 64.525 52.787 67.095 52.843 ;
      RECT 64.571 52.741 67.141 52.797 ;
      RECT 64.617 52.695 67.187 52.751 ;
      RECT 64.663 52.649 67.233 52.705 ;
      RECT 64.709 52.603 67.279 52.659 ;
      RECT 64.755 52.557 67.325 52.613 ;
      RECT 64.801 52.511 67.371 52.567 ;
      RECT 64.847 52.465 67.417 52.521 ;
      RECT 64.893 52.419 67.463 52.475 ;
      RECT 64.939 52.373 67.509 52.429 ;
      RECT 64.985 52.327 67.555 52.383 ;
      RECT 65.031 52.281 67.601 52.337 ;
      RECT 65.077 52.235 67.647 52.291 ;
      RECT 65.123 52.189 67.693 52.245 ;
      RECT 65.169 52.143 67.739 52.199 ;
      RECT 65.215 52.097 67.785 52.153 ;
      RECT 65.261 52.051 67.831 52.107 ;
      RECT 65.307 52.005 67.877 52.061 ;
      RECT 65.353 51.959 67.923 52.015 ;
      RECT 65.399 51.913 67.969 51.969 ;
      RECT 65.445 51.867 68.015 51.923 ;
      RECT 65.491 51.821 68.061 51.877 ;
      RECT 65.537 51.775 68.107 51.831 ;
      RECT 65.583 51.729 68.153 51.785 ;
      RECT 65.629 51.683 68.199 51.739 ;
      RECT 65.675 51.637 68.245 51.693 ;
      RECT 65.721 51.591 68.291 51.647 ;
      RECT 65.767 51.545 68.337 51.601 ;
      RECT 65.813 51.499 68.383 51.555 ;
      RECT 65.859 51.453 68.429 51.509 ;
      RECT 65.905 51.407 68.475 51.463 ;
      RECT 65.951 51.361 68.521 51.417 ;
      RECT 65.997 51.315 68.567 51.371 ;
      RECT 66.043 51.269 68.613 51.325 ;
      RECT 66.089 51.223 68.659 51.279 ;
      RECT 66.135 51.177 68.705 51.233 ;
      RECT 66.181 51.131 68.751 51.187 ;
      RECT 66.227 51.085 68.797 51.141 ;
      RECT 66.273 51.039 68.843 51.095 ;
      RECT 66.319 50.993 68.889 51.049 ;
      RECT 66.365 50.947 68.935 51.003 ;
      RECT 66.411 50.901 68.981 50.957 ;
      RECT 66.457 50.855 69.027 50.911 ;
      RECT 66.503 50.809 69.073 50.865 ;
      RECT 66.549 50.763 69.119 50.819 ;
      RECT 66.595 50.717 69.165 50.773 ;
      RECT 66.641 50.671 69.211 50.727 ;
      RECT 66.687 50.625 69.257 50.681 ;
      RECT 66.733 50.579 69.303 50.635 ;
      RECT 66.779 50.533 69.349 50.589 ;
      RECT 66.825 50.487 69.395 50.543 ;
      RECT 66.871 50.441 69.441 50.497 ;
      RECT 66.917 50.395 69.487 50.451 ;
      RECT 66.963 50.349 69.533 50.405 ;
      RECT 67.009 50.303 69.579 50.359 ;
      RECT 67.055 50.257 69.625 50.313 ;
      RECT 67.101 50.211 69.671 50.267 ;
      RECT 67.147 50.165 69.717 50.221 ;
      RECT 69.677 47.652 69.717 50.221 ;
      RECT 67.193 50.119 69.763 50.175 ;
      RECT 69.69 47.622 69.763 50.175 ;
      RECT 67.239 50.073 69.809 50.129 ;
      RECT 69.736 47.576 69.809 50.129 ;
      RECT 67.285 50.027 69.855 50.083 ;
      RECT 69.782 47.53 69.855 50.083 ;
      RECT 67.331 49.981 69.901 50.037 ;
      RECT 69.828 47.484 69.901 50.037 ;
      RECT 67.377 49.935 69.947 49.991 ;
      RECT 69.874 47.438 69.947 49.991 ;
      RECT 67.423 49.889 69.993 49.945 ;
      RECT 69.92 47.392 69.993 49.945 ;
      RECT 67.469 49.843 70.039 49.899 ;
      RECT 69.966 47.346 70.039 49.899 ;
      RECT 67.515 49.797 70.085 49.853 ;
      RECT 70.012 47.3 70.085 49.853 ;
      RECT 67.561 49.751 70.131 49.807 ;
      RECT 70.058 47.254 70.131 49.807 ;
      RECT 67.607 49.705 70.177 49.761 ;
      RECT 70.104 47.208 70.177 49.761 ;
      RECT 67.653 49.659 70.223 49.715 ;
      RECT 70.15 47.162 70.223 49.715 ;
      RECT 67.699 49.613 70.269 49.669 ;
      RECT 70.196 47.116 70.269 49.669 ;
      RECT 67.745 49.567 70.315 49.623 ;
      RECT 70.242 47.07 70.315 49.623 ;
      RECT 67.791 49.521 70.361 49.577 ;
      RECT 70.288 47.024 70.361 49.577 ;
      RECT 67.837 49.475 70.407 49.531 ;
      RECT 70.334 46.978 70.407 49.531 ;
      RECT 67.883 49.429 70.453 49.485 ;
      RECT 70.38 46.932 70.453 49.485 ;
      RECT 67.929 49.383 70.499 49.439 ;
      RECT 70.426 46.886 70.499 49.439 ;
      RECT 67.975 49.337 70.545 49.393 ;
      RECT 70.472 46.84 70.545 49.393 ;
      RECT 68.021 49.291 70.591 49.347 ;
      RECT 70.518 46.794 70.591 49.347 ;
      RECT 68.067 49.245 70.637 49.301 ;
      RECT 70.564 46.748 70.637 49.301 ;
      RECT 68.113 49.199 70.683 49.255 ;
      RECT 70.61 46.702 70.683 49.255 ;
      RECT 68.159 49.153 70.729 49.209 ;
      RECT 70.656 46.656 70.729 49.209 ;
      RECT 68.205 49.107 70.775 49.163 ;
      RECT 70.702 46.61 70.775 49.163 ;
      RECT 68.251 49.061 70.821 49.117 ;
      RECT 70.748 46.564 70.821 49.117 ;
      RECT 68.297 49.015 70.867 49.071 ;
      RECT 70.794 46.518 70.867 49.071 ;
      RECT 68.343 48.969 70.913 49.025 ;
      RECT 70.84 46.472 70.913 49.025 ;
      RECT 68.389 48.923 70.959 48.979 ;
      RECT 70.886 46.426 70.959 48.979 ;
      RECT 68.435 48.877 71.005 48.933 ;
      RECT 70.932 46.38 71.005 48.933 ;
      RECT 68.481 48.831 71.051 48.887 ;
      RECT 70.978 46.334 71.051 48.887 ;
      RECT 68.527 48.785 71.097 48.841 ;
      RECT 71.024 46.288 71.097 48.841 ;
      RECT 68.573 48.739 71.143 48.795 ;
      RECT 71.07 46.242 71.143 48.795 ;
      RECT 68.619 48.693 71.189 48.749 ;
      RECT 71.116 46.196 71.189 48.749 ;
      RECT 68.665 48.647 71.235 48.703 ;
      RECT 71.162 46.15 71.235 48.703 ;
      RECT 68.711 48.601 71.281 48.657 ;
      RECT 71.208 46.104 71.281 48.657 ;
      RECT 68.757 48.555 71.327 48.611 ;
      RECT 71.254 46.058 71.327 48.611 ;
      RECT 68.803 48.509 71.373 48.565 ;
      RECT 71.3 46.012 71.373 48.565 ;
      RECT 68.849 48.463 71.419 48.519 ;
      RECT 71.346 45.966 71.419 48.519 ;
      RECT 68.895 48.417 71.465 48.473 ;
      RECT 71.392 45.92 71.465 48.473 ;
      RECT 68.941 48.371 71.511 48.427 ;
      RECT 71.438 45.874 71.511 48.427 ;
      RECT 68.987 48.325 71.557 48.381 ;
      RECT 71.484 45.828 71.557 48.381 ;
      RECT 69.033 48.279 71.603 48.335 ;
      RECT 71.53 45.782 71.603 48.335 ;
      RECT 69.079 48.233 71.649 48.289 ;
      RECT 71.576 45.736 71.649 48.289 ;
      RECT 69.125 48.187 71.695 48.243 ;
      RECT 71.622 45.69 71.695 48.243 ;
      RECT 69.171 48.141 71.741 48.197 ;
      RECT 71.668 45.644 71.741 48.197 ;
      RECT 69.217 48.095 71.787 48.151 ;
      RECT 71.714 45.598 71.787 48.151 ;
      RECT 69.263 48.049 71.833 48.105 ;
      RECT 71.76 45.552 71.833 48.105 ;
      RECT 69.309 48.003 71.879 48.059 ;
      RECT 71.806 45.506 71.879 48.059 ;
      RECT 69.355 47.957 71.925 48.013 ;
      RECT 71.852 45.46 71.925 48.013 ;
      RECT 69.401 47.911 71.971 47.967 ;
      RECT 71.898 45.414 71.971 47.967 ;
      RECT 69.447 47.865 72.017 47.921 ;
      RECT 71.944 45.368 72.017 47.921 ;
      RECT 69.493 47.819 72.063 47.875 ;
      RECT 71.99 45.322 72.063 47.875 ;
      RECT 69.539 47.773 72.109 47.829 ;
      RECT 72.036 45.276 72.109 47.829 ;
      RECT 69.585 47.727 72.155 47.783 ;
      RECT 72.082 45.23 72.155 47.783 ;
      RECT 69.631 47.681 72.201 47.737 ;
      RECT 72.128 45.184 72.201 47.737 ;
      RECT 72.174 45.138 72.247 47.691 ;
      RECT 72.22 45.092 72.293 47.645 ;
      RECT 72.266 45.046 72.339 47.599 ;
      RECT 72.312 45 72.385 47.553 ;
      RECT 72.358 44.954 72.431 47.507 ;
      RECT 72.404 44.908 72.477 47.461 ;
      RECT 72.45 44.862 72.523 47.415 ;
      RECT 72.496 44.816 72.569 47.369 ;
      RECT 72.542 44.77 72.615 47.323 ;
      RECT 72.588 44.724 72.661 47.277 ;
      RECT 72.634 44.678 72.707 47.231 ;
      RECT 72.68 44.632 72.753 47.185 ;
      RECT 72.726 44.586 72.799 47.139 ;
      RECT 72.772 44.54 72.845 47.093 ;
      RECT 72.818 44.494 72.891 47.047 ;
      RECT 72.864 44.448 72.937 47.001 ;
      RECT 72.91 44.402 72.983 46.955 ;
      RECT 72.956 44.356 73.029 46.909 ;
      RECT 73.002 44.31 73.075 46.863 ;
      RECT 73.048 44.264 73.121 46.817 ;
      RECT 73.094 44.218 73.167 46.771 ;
      RECT 73.14 44.172 73.213 46.725 ;
      RECT 73.186 44.126 73.259 46.679 ;
      RECT 73.232 44.08 73.305 46.633 ;
      RECT 73.278 44.034 73.351 46.587 ;
      RECT 73.324 43.988 73.397 46.541 ;
      RECT 73.37 43.942 73.443 46.495 ;
      RECT 73.416 43.896 73.489 46.449 ;
      RECT 73.462 43.85 73.535 46.403 ;
      RECT 73.508 43.804 73.581 46.357 ;
      RECT 73.554 43.758 73.627 46.311 ;
      RECT 73.6 43.712 73.673 46.265 ;
      RECT 73.646 43.666 73.719 46.219 ;
      RECT 73.692 43.62 73.765 46.173 ;
      RECT 73.738 43.574 73.811 46.127 ;
      RECT 73.784 43.528 73.857 46.081 ;
      RECT 73.83 43.482 73.903 46.035 ;
      RECT 73.876 43.436 73.949 45.989 ;
      RECT 73.922 43.39 73.995 45.943 ;
      RECT 73.968 43.344 74.041 45.897 ;
      RECT 74.014 43.298 74.087 45.851 ;
      RECT 74.06 43.252 74.133 45.805 ;
      RECT 74.106 43.206 74.179 45.759 ;
      RECT 74.152 43.16 74.225 45.713 ;
      RECT 74.198 43.114 74.271 45.667 ;
      RECT 74.244 43.068 74.317 45.621 ;
      RECT 74.29 43.022 74.363 45.575 ;
      RECT 74.336 42.976 74.409 45.529 ;
      RECT 74.382 42.93 74.455 45.483 ;
      RECT 74.428 42.884 74.501 45.437 ;
      RECT 74.474 42.838 74.547 45.391 ;
      RECT 74.52 42.792 74.593 45.345 ;
      RECT 74.566 42.746 74.639 45.299 ;
      RECT 74.612 42.699 74.685 45.253 ;
      RECT 74.658 42.675 74.731 45.207 ;
      RECT 74.658 42.675 74.777 45.161 ;
      RECT 74.658 42.675 74.823 45.115 ;
      RECT 74.658 42.675 74.869 45.069 ;
      RECT 74.658 42.675 74.915 45.023 ;
      RECT 74.658 42.675 74.961 44.977 ;
      RECT 74.658 42.675 75.007 44.931 ;
      RECT 74.658 42.675 75.053 44.885 ;
      RECT 74.658 42.675 75.099 44.839 ;
      RECT 74.658 42.675 75.145 44.793 ;
      RECT 74.658 42.675 75.191 44.747 ;
      RECT 74.658 42.675 75.237 44.701 ;
      RECT 74.658 42.675 75.283 44.655 ;
      RECT 74.658 42.675 75.329 44.609 ;
      RECT 74.658 42.675 75.375 44.563 ;
      RECT 74.658 42.675 75.421 44.517 ;
      RECT 74.658 42.675 75.467 44.471 ;
      RECT 74.658 42.675 75.513 44.425 ;
      RECT 74.658 42.675 75.559 44.379 ;
      RECT 74.658 42.675 75.605 44.333 ;
      RECT 74.658 42.675 75.651 44.287 ;
      RECT 74.658 42.675 75.697 44.241 ;
      RECT 74.658 42.675 75.743 44.195 ;
      RECT 74.658 42.675 75.789 44.149 ;
      RECT 74.658 42.675 75.835 44.103 ;
      RECT 74.658 42.675 75.881 44.057 ;
      RECT 74.658 42.675 75.927 44.011 ;
      RECT 74.658 42.675 75.973 43.965 ;
      RECT 74.658 42.675 76.019 43.919 ;
      RECT 74.658 42.675 76.065 43.873 ;
      RECT 73.508 43.804 76.09 43.837 ;
      RECT 74.658 42.675 110 43.825 ;
      RECT 56.175 81.387 57.325 110 ;
      RECT 56.175 81.387 57.371 82.562 ;
      RECT 56.175 81.387 57.417 82.516 ;
      RECT 56.175 81.387 57.463 82.47 ;
      RECT 56.175 81.387 57.509 82.424 ;
      RECT 56.175 81.387 57.555 82.378 ;
      RECT 56.175 81.387 57.601 82.332 ;
      RECT 56.175 81.387 57.647 82.286 ;
      RECT 56.175 81.387 57.693 82.24 ;
      RECT 56.175 81.387 57.739 82.194 ;
      RECT 56.175 81.387 57.785 82.148 ;
      RECT 56.175 81.387 57.831 82.102 ;
      RECT 56.175 81.387 57.877 82.056 ;
      RECT 56.175 81.387 57.923 82.01 ;
      RECT 56.175 81.387 57.969 81.964 ;
      RECT 56.175 81.387 58.015 81.918 ;
      RECT 56.175 81.387 58.061 81.872 ;
      RECT 56.175 81.387 58.107 81.826 ;
      RECT 56.175 81.387 58.153 81.78 ;
      RECT 56.175 81.387 58.199 81.734 ;
      RECT 56.175 81.387 58.245 81.688 ;
      RECT 56.175 81.387 58.291 81.642 ;
      RECT 56.175 81.387 58.337 81.596 ;
      RECT 56.175 81.387 58.383 81.55 ;
      RECT 56.175 81.387 58.429 81.504 ;
      RECT 56.175 81.387 58.475 81.458 ;
      RECT 56.221 81.341 58.521 81.412 ;
      RECT 56.267 81.295 58.567 81.366 ;
      RECT 56.313 81.249 58.613 81.32 ;
      RECT 56.359 81.203 58.659 81.274 ;
      RECT 56.405 81.157 58.705 81.228 ;
      RECT 56.451 81.111 58.751 81.182 ;
      RECT 56.497 81.065 58.797 81.136 ;
      RECT 56.543 81.019 58.843 81.09 ;
      RECT 56.589 80.973 58.889 81.044 ;
      RECT 56.635 80.927 58.935 80.998 ;
      RECT 56.681 80.881 58.981 80.952 ;
      RECT 56.727 80.835 59.027 80.906 ;
      RECT 56.773 80.789 59.073 80.86 ;
      RECT 56.819 80.743 59.119 80.814 ;
      RECT 56.865 80.697 59.165 80.768 ;
      RECT 56.911 80.651 59.211 80.722 ;
      RECT 56.957 80.605 59.257 80.676 ;
      RECT 57.003 80.559 59.303 80.63 ;
      RECT 57.049 80.513 59.349 80.584 ;
      RECT 57.095 80.467 59.395 80.538 ;
      RECT 57.141 80.421 59.441 80.492 ;
      RECT 57.187 80.375 59.487 80.446 ;
      RECT 57.233 80.329 59.533 80.4 ;
      RECT 57.279 80.283 59.579 80.354 ;
      RECT 57.325 80.237 59.625 80.308 ;
      RECT 57.371 80.191 59.671 80.262 ;
      RECT 57.417 80.145 59.717 80.216 ;
      RECT 57.463 80.099 59.763 80.17 ;
      RECT 57.509 80.053 59.809 80.124 ;
      RECT 57.555 80.007 59.855 80.078 ;
      RECT 57.601 79.961 59.901 80.032 ;
      RECT 57.647 79.915 59.947 79.986 ;
      RECT 57.693 79.869 59.993 79.94 ;
      RECT 57.739 79.823 60.039 79.894 ;
      RECT 57.785 79.777 60.085 79.848 ;
      RECT 57.831 79.731 60.131 79.802 ;
      RECT 57.877 79.685 60.177 79.756 ;
      RECT 57.923 79.639 60.223 79.71 ;
      RECT 57.969 79.593 60.269 79.664 ;
      RECT 58.015 79.547 60.315 79.618 ;
      RECT 58.061 79.501 60.361 79.572 ;
      RECT 58.107 79.455 60.407 79.526 ;
      RECT 58.153 79.409 60.453 79.48 ;
      RECT 58.199 79.363 60.499 79.434 ;
      RECT 58.245 79.317 60.545 79.388 ;
      RECT 58.291 79.271 60.591 79.342 ;
      RECT 58.337 79.225 60.637 79.296 ;
      RECT 58.383 79.179 60.683 79.25 ;
      RECT 58.429 79.133 60.729 79.204 ;
      RECT 58.475 79.087 60.775 79.158 ;
      RECT 58.521 79.041 60.821 79.112 ;
      RECT 58.567 78.995 60.867 79.066 ;
      RECT 58.613 78.949 60.913 79.02 ;
      RECT 58.659 78.903 60.959 78.974 ;
      RECT 58.705 78.857 61.005 78.928 ;
      RECT 58.751 78.811 61.051 78.882 ;
      RECT 58.797 78.765 61.097 78.836 ;
      RECT 58.843 78.719 61.143 78.79 ;
      RECT 58.889 78.673 61.189 78.744 ;
      RECT 58.935 78.627 61.235 78.698 ;
      RECT 58.981 78.581 61.281 78.652 ;
      RECT 59.027 78.535 61.327 78.606 ;
      RECT 59.073 78.489 61.373 78.56 ;
      RECT 59.119 78.443 61.419 78.514 ;
      RECT 59.165 78.397 61.465 78.468 ;
      RECT 59.211 78.351 61.511 78.422 ;
      RECT 59.257 78.305 61.557 78.376 ;
      RECT 59.303 78.259 61.603 78.33 ;
      RECT 59.349 78.213 61.649 78.284 ;
      RECT 59.395 78.167 61.695 78.238 ;
      RECT 59.441 78.121 61.741 78.192 ;
      RECT 59.487 78.075 61.787 78.146 ;
      RECT 59.533 78.029 61.833 78.1 ;
      RECT 59.579 77.983 61.879 78.054 ;
      RECT 59.625 77.937 61.925 78.008 ;
      RECT 59.671 77.891 61.971 77.962 ;
      RECT 59.717 77.845 62.017 77.916 ;
      RECT 59.763 77.799 62.063 77.87 ;
      RECT 59.809 77.753 62.109 77.824 ;
      RECT 59.855 77.707 62.155 77.778 ;
      RECT 59.901 77.661 62.201 77.732 ;
      RECT 59.947 77.615 62.247 77.686 ;
      RECT 59.993 77.569 62.293 77.64 ;
      RECT 60.039 77.523 62.339 77.594 ;
      RECT 60.085 77.477 62.385 77.548 ;
      RECT 60.131 77.431 62.431 77.502 ;
      RECT 60.177 77.385 62.477 77.456 ;
      RECT 60.223 77.339 62.523 77.41 ;
      RECT 60.269 77.293 62.569 77.364 ;
      RECT 60.315 77.247 62.615 77.318 ;
      RECT 60.361 77.201 62.661 77.272 ;
      RECT 60.407 77.155 62.707 77.226 ;
      RECT 60.453 77.109 62.753 77.18 ;
      RECT 60.499 77.063 62.799 77.134 ;
      RECT 60.545 77.017 62.845 77.088 ;
      RECT 60.591 76.971 62.891 77.042 ;
      RECT 60.637 76.925 62.937 76.996 ;
      RECT 60.683 76.879 62.983 76.95 ;
      RECT 60.729 76.833 63.029 76.904 ;
      RECT 60.775 76.787 63.075 76.858 ;
      RECT 60.821 76.741 63.121 76.812 ;
      RECT 60.867 76.695 63.167 76.766 ;
      RECT 60.913 76.649 63.213 76.72 ;
      RECT 60.959 76.603 63.259 76.674 ;
      RECT 61.005 76.557 63.305 76.628 ;
      RECT 61.005 76.557 63.325 76.595 ;
      RECT 61.051 76.511 63.371 76.562 ;
      RECT 63.305 74.257 63.371 76.562 ;
      RECT 61.097 76.465 63.417 76.516 ;
      RECT 63.351 74.211 63.417 76.516 ;
      RECT 61.143 76.419 63.463 76.47 ;
      RECT 63.397 74.165 63.463 76.47 ;
      RECT 61.189 76.373 63.509 76.424 ;
      RECT 63.443 74.119 63.509 76.424 ;
      RECT 61.235 76.327 63.555 76.378 ;
      RECT 63.489 74.073 63.555 76.378 ;
      RECT 61.281 76.281 63.601 76.332 ;
      RECT 63.535 74.027 63.601 76.332 ;
      RECT 61.327 76.235 63.647 76.286 ;
      RECT 63.581 73.981 63.647 76.286 ;
      RECT 61.373 76.189 63.693 76.24 ;
      RECT 63.627 73.935 63.693 76.24 ;
      RECT 61.419 76.143 63.739 76.194 ;
      RECT 63.673 73.889 63.739 76.194 ;
      RECT 61.465 76.097 63.785 76.148 ;
      RECT 63.719 73.843 63.785 76.148 ;
      RECT 61.511 76.051 63.831 76.102 ;
      RECT 63.765 73.797 63.831 76.102 ;
      RECT 61.557 76.005 63.877 76.056 ;
      RECT 63.811 73.751 63.877 76.056 ;
      RECT 61.603 75.959 63.923 76.01 ;
      RECT 63.857 73.705 63.923 76.01 ;
      RECT 61.649 75.913 63.969 75.964 ;
      RECT 63.903 73.659 63.969 75.964 ;
      RECT 61.695 75.867 64.015 75.918 ;
      RECT 63.949 73.613 64.015 75.918 ;
      RECT 61.741 75.821 64.061 75.872 ;
      RECT 63.995 73.567 64.061 75.872 ;
      RECT 61.787 75.775 64.107 75.826 ;
      RECT 64.041 73.521 64.107 75.826 ;
      RECT 61.833 75.729 64.153 75.78 ;
      RECT 64.087 73.475 64.153 75.78 ;
      RECT 61.879 75.683 64.199 75.734 ;
      RECT 64.133 73.429 64.199 75.734 ;
      RECT 61.925 75.637 64.245 75.688 ;
      RECT 64.179 73.383 64.245 75.688 ;
      RECT 61.971 75.591 64.291 75.642 ;
      RECT 64.225 73.337 64.291 75.642 ;
      RECT 62.017 75.545 64.337 75.596 ;
      RECT 64.271 73.291 64.337 75.596 ;
      RECT 62.063 75.499 64.383 75.55 ;
      RECT 64.317 73.245 64.383 75.55 ;
      RECT 62.109 75.453 64.429 75.504 ;
      RECT 64.363 73.199 64.429 75.504 ;
      RECT 62.155 75.407 64.475 75.458 ;
      RECT 64.409 73.153 64.475 75.458 ;
      RECT 62.201 75.361 64.521 75.412 ;
      RECT 64.455 73.107 64.521 75.412 ;
      RECT 62.247 75.315 64.567 75.366 ;
      RECT 64.501 73.061 64.567 75.366 ;
      RECT 62.293 75.269 64.613 75.32 ;
      RECT 64.547 73.015 64.613 75.32 ;
      RECT 62.339 75.223 64.659 75.274 ;
      RECT 64.593 72.969 64.659 75.274 ;
      RECT 62.385 75.177 64.705 75.228 ;
      RECT 64.639 72.923 64.705 75.228 ;
      RECT 62.431 75.131 64.751 75.182 ;
      RECT 64.685 72.877 64.751 75.182 ;
      RECT 62.477 75.085 64.797 75.136 ;
      RECT 64.731 72.831 64.797 75.136 ;
      RECT 62.523 75.039 64.843 75.09 ;
      RECT 64.777 72.785 64.843 75.09 ;
      RECT 62.569 74.993 64.889 75.044 ;
      RECT 64.823 72.739 64.889 75.044 ;
      RECT 62.615 74.947 64.935 74.998 ;
      RECT 64.869 72.693 64.935 74.998 ;
      RECT 62.661 74.901 64.981 74.952 ;
      RECT 64.915 72.647 64.981 74.952 ;
      RECT 62.707 74.855 65.027 74.906 ;
      RECT 64.961 72.601 65.027 74.906 ;
      RECT 62.753 74.809 65.073 74.86 ;
      RECT 65.007 72.555 65.073 74.86 ;
      RECT 62.799 74.763 65.119 74.814 ;
      RECT 65.053 72.509 65.119 74.814 ;
      RECT 62.845 74.717 65.165 74.768 ;
      RECT 65.099 72.463 65.165 74.768 ;
      RECT 62.891 74.671 65.211 74.722 ;
      RECT 65.145 72.417 65.211 74.722 ;
      RECT 62.937 74.625 65.257 74.676 ;
      RECT 65.191 72.371 65.257 74.676 ;
      RECT 62.983 74.579 65.303 74.63 ;
      RECT 65.237 72.325 65.303 74.63 ;
      RECT 63.029 74.533 65.349 74.584 ;
      RECT 65.283 72.279 65.349 74.584 ;
      RECT 63.075 74.487 65.395 74.538 ;
      RECT 65.329 72.233 65.395 74.538 ;
      RECT 63.121 74.441 65.441 74.492 ;
      RECT 65.375 72.187 65.441 74.492 ;
      RECT 63.167 74.395 65.487 74.446 ;
      RECT 65.421 72.141 65.487 74.446 ;
      RECT 63.213 74.349 65.533 74.4 ;
      RECT 65.467 72.095 65.533 74.4 ;
      RECT 63.259 74.303 65.579 74.354 ;
      RECT 65.513 72.049 65.579 74.354 ;
      RECT 65.559 72.003 65.625 74.308 ;
      RECT 65.605 71.957 65.671 74.262 ;
      RECT 65.651 71.911 65.717 74.216 ;
      RECT 65.697 71.865 65.763 74.17 ;
      RECT 65.743 71.819 65.809 74.124 ;
      RECT 65.789 71.773 65.855 74.078 ;
      RECT 65.835 71.727 65.901 74.032 ;
      RECT 65.881 71.681 65.947 73.986 ;
      RECT 65.927 71.635 65.993 73.94 ;
      RECT 65.973 71.589 66.039 73.894 ;
      RECT 66.019 71.543 66.085 73.848 ;
      RECT 66.065 71.497 66.131 73.802 ;
      RECT 66.111 71.451 66.177 73.756 ;
      RECT 66.157 71.405 66.223 73.71 ;
      RECT 66.203 71.359 66.269 73.664 ;
      RECT 66.249 71.313 66.315 73.618 ;
      RECT 66.295 71.267 66.361 73.572 ;
      RECT 66.341 71.221 66.407 73.526 ;
      RECT 66.387 71.175 66.453 73.48 ;
      RECT 66.433 71.129 66.499 73.434 ;
      RECT 66.479 71.083 66.545 73.388 ;
      RECT 66.525 71.037 66.591 73.342 ;
      RECT 66.571 70.991 66.637 73.296 ;
      RECT 66.617 70.945 66.683 73.25 ;
      RECT 66.663 70.899 66.729 73.204 ;
      RECT 66.709 70.853 66.775 73.158 ;
      RECT 66.755 70.807 66.821 73.112 ;
      RECT 66.801 70.761 66.867 73.066 ;
      RECT 66.847 70.715 66.913 73.02 ;
      RECT 66.893 70.669 66.959 72.974 ;
      RECT 66.939 70.623 67.005 72.928 ;
      RECT 66.985 70.577 67.051 72.882 ;
      RECT 67.031 70.531 67.097 72.836 ;
      RECT 67.077 70.485 67.143 72.79 ;
      RECT 67.123 70.439 67.189 72.744 ;
      RECT 67.169 70.393 67.235 72.698 ;
      RECT 67.215 70.347 67.281 72.652 ;
      RECT 67.261 70.301 67.327 72.606 ;
      RECT 67.307 70.255 67.373 72.56 ;
      RECT 67.353 70.209 67.419 72.514 ;
      RECT 67.399 70.163 67.465 72.468 ;
      RECT 67.445 70.117 67.511 72.422 ;
      RECT 67.491 70.071 67.557 72.376 ;
      RECT 67.537 70.025 67.603 72.33 ;
      RECT 67.583 69.979 67.649 72.284 ;
      RECT 67.629 69.933 67.695 72.238 ;
      RECT 67.675 69.887 67.741 72.192 ;
      RECT 67.721 69.841 67.787 72.146 ;
      RECT 67.767 69.795 67.833 72.1 ;
      RECT 67.813 69.749 67.879 72.054 ;
      RECT 67.859 69.703 67.925 72.008 ;
      RECT 67.905 69.657 67.971 71.962 ;
      RECT 67.951 69.611 68.017 71.916 ;
      RECT 67.997 69.565 68.063 71.87 ;
      RECT 68.043 69.519 68.109 71.824 ;
      RECT 68.089 69.473 68.155 71.778 ;
      RECT 68.135 69.427 68.201 71.732 ;
      RECT 68.181 69.381 68.247 71.686 ;
      RECT 68.227 69.335 68.293 71.64 ;
      RECT 68.273 69.289 68.339 71.594 ;
      RECT 68.319 69.243 68.385 71.548 ;
      RECT 68.365 69.197 68.431 71.502 ;
      RECT 68.411 69.151 68.477 71.456 ;
      RECT 68.457 69.105 68.523 71.41 ;
      RECT 68.503 69.059 68.569 71.364 ;
      RECT 68.549 69.013 68.615 71.318 ;
      RECT 68.595 68.967 68.661 71.272 ;
      RECT 68.641 68.921 68.707 71.226 ;
      RECT 68.687 68.875 68.753 71.18 ;
      RECT 68.733 68.829 68.799 71.134 ;
      RECT 68.779 68.783 68.845 71.088 ;
      RECT 68.825 68.737 68.891 71.042 ;
      RECT 68.871 68.691 68.937 70.996 ;
      RECT 68.917 68.645 68.983 70.95 ;
      RECT 68.963 68.599 69.029 70.904 ;
      RECT 69.009 68.553 69.075 70.858 ;
      RECT 69.055 68.507 69.121 70.812 ;
      RECT 69.101 68.461 69.167 70.766 ;
      RECT 69.147 68.415 69.213 70.72 ;
      RECT 69.193 68.369 69.259 70.674 ;
      RECT 69.239 68.323 69.305 70.628 ;
      RECT 69.285 68.277 69.351 70.582 ;
      RECT 69.331 68.231 69.397 70.536 ;
      RECT 69.377 68.185 69.443 70.49 ;
      RECT 69.423 68.139 69.489 70.444 ;
      RECT 69.469 68.093 69.535 70.398 ;
      RECT 69.515 68.047 69.581 70.352 ;
      RECT 69.561 68.001 69.627 70.306 ;
      RECT 69.607 67.955 69.673 70.26 ;
      RECT 69.653 67.909 69.719 70.214 ;
      RECT 69.699 67.863 69.765 70.168 ;
      RECT 69.745 67.817 69.811 70.122 ;
      RECT 69.791 67.771 69.857 70.076 ;
      RECT 69.837 67.725 69.903 70.03 ;
      RECT 69.883 67.679 69.949 69.984 ;
      RECT 69.929 67.633 69.995 69.938 ;
      RECT 69.975 67.587 70.041 69.892 ;
      RECT 70.021 67.541 70.087 69.846 ;
      RECT 70.067 67.495 70.133 69.8 ;
      RECT 70.113 67.449 70.179 69.754 ;
      RECT 70.159 67.403 70.225 69.708 ;
      RECT 70.205 67.357 70.271 69.662 ;
      RECT 70.251 67.311 70.317 69.616 ;
      RECT 70.297 67.265 70.363 69.57 ;
      RECT 70.343 67.219 70.409 69.524 ;
      RECT 70.389 67.173 70.455 69.478 ;
      RECT 70.435 67.127 70.501 69.432 ;
      RECT 70.481 67.081 70.547 69.386 ;
      RECT 70.527 67.035 70.593 69.34 ;
      RECT 70.573 66.989 70.639 69.294 ;
      RECT 70.619 66.943 70.685 69.248 ;
      RECT 70.665 66.897 70.731 69.202 ;
      RECT 70.711 66.851 70.777 69.156 ;
      RECT 70.757 66.805 70.823 69.11 ;
      RECT 70.803 66.759 70.869 69.064 ;
      RECT 70.849 66.713 70.915 69.018 ;
      RECT 70.895 66.667 70.961 68.972 ;
      RECT 70.941 66.621 71.007 68.926 ;
      RECT 70.987 66.575 71.053 68.88 ;
      RECT 71.033 66.529 71.099 68.834 ;
      RECT 71.079 66.483 71.145 68.788 ;
      RECT 71.125 66.437 71.191 68.742 ;
      RECT 71.171 66.391 71.237 68.696 ;
      RECT 71.217 66.345 71.283 68.65 ;
      RECT 71.263 66.299 71.329 68.604 ;
      RECT 71.309 66.253 71.375 68.558 ;
      RECT 71.355 66.207 71.421 68.512 ;
      RECT 71.401 66.161 71.467 68.466 ;
      RECT 71.447 66.115 71.513 68.42 ;
      RECT 71.493 66.069 71.559 68.374 ;
      RECT 71.539 66.023 71.605 68.328 ;
      RECT 71.585 65.977 71.651 68.282 ;
      RECT 71.631 65.931 71.697 68.236 ;
      RECT 71.677 65.885 71.743 68.19 ;
      RECT 71.723 65.839 71.789 68.144 ;
      RECT 71.769 65.793 71.835 68.098 ;
      RECT 71.815 65.747 71.881 68.052 ;
      RECT 71.861 65.701 71.927 68.006 ;
      RECT 71.907 65.655 71.973 67.96 ;
      RECT 71.953 65.609 72.019 67.914 ;
      RECT 71.999 65.563 72.065 67.868 ;
      RECT 72.045 65.517 72.111 67.822 ;
      RECT 72.091 65.471 72.157 67.776 ;
      RECT 72.137 65.425 72.203 67.73 ;
      RECT 72.183 65.379 72.249 67.684 ;
      RECT 72.229 65.333 72.295 67.638 ;
      RECT 72.275 65.287 72.341 67.592 ;
      RECT 72.321 65.241 72.387 67.546 ;
      RECT 72.367 65.195 72.433 67.5 ;
      RECT 72.413 65.149 72.479 67.454 ;
      RECT 72.459 65.103 72.525 67.408 ;
      RECT 72.505 65.057 72.571 67.362 ;
      RECT 72.551 65.011 72.617 67.316 ;
      RECT 72.597 64.965 72.663 67.27 ;
      RECT 72.643 64.919 72.709 67.224 ;
      RECT 72.689 64.873 72.755 67.178 ;
      RECT 72.735 64.827 72.801 67.132 ;
      RECT 72.781 64.781 72.847 67.086 ;
      RECT 72.827 64.735 72.893 67.04 ;
      RECT 72.873 64.689 72.939 66.994 ;
      RECT 72.919 64.643 72.985 66.948 ;
      RECT 72.965 64.597 73.031 66.902 ;
      RECT 73.011 64.551 73.077 66.856 ;
      RECT 73.057 64.505 73.123 66.81 ;
      RECT 73.103 64.459 73.169 66.764 ;
      RECT 73.149 64.413 73.215 66.718 ;
      RECT 73.195 64.367 73.261 66.672 ;
      RECT 73.241 64.321 73.307 66.626 ;
      RECT 73.287 64.275 73.353 66.58 ;
      RECT 73.333 64.229 73.399 66.534 ;
      RECT 73.379 64.183 73.445 66.488 ;
      RECT 73.425 64.137 73.491 66.442 ;
      RECT 73.471 64.091 73.537 66.396 ;
      RECT 73.517 64.045 73.583 66.35 ;
      RECT 73.563 63.999 73.629 66.304 ;
      RECT 73.609 63.953 73.675 66.258 ;
      RECT 73.655 63.907 73.721 66.212 ;
      RECT 73.701 63.861 73.767 66.166 ;
      RECT 73.747 63.815 73.813 66.12 ;
      RECT 73.793 63.769 73.859 66.074 ;
      RECT 73.839 63.723 73.905 66.028 ;
      RECT 73.885 63.677 73.951 65.982 ;
      RECT 73.931 63.631 73.997 65.936 ;
      RECT 73.977 63.585 74.043 65.89 ;
      RECT 74.023 63.539 74.089 65.844 ;
      RECT 74.069 63.493 74.135 65.798 ;
      RECT 74.115 63.447 74.181 65.752 ;
      RECT 74.161 63.401 74.227 65.706 ;
      RECT 74.207 63.355 74.273 65.66 ;
      RECT 74.253 63.309 74.319 65.614 ;
      RECT 74.299 63.263 74.365 65.568 ;
      RECT 74.345 63.217 74.411 65.522 ;
      RECT 74.391 63.171 74.457 65.476 ;
      RECT 74.437 63.125 74.503 65.43 ;
      RECT 74.483 63.079 74.549 65.384 ;
      RECT 74.529 63.033 74.595 65.338 ;
      RECT 74.575 62.987 74.641 65.292 ;
      RECT 74.621 62.941 74.687 65.246 ;
      RECT 74.667 62.895 74.733 65.2 ;
      RECT 74.713 62.849 74.779 65.154 ;
      RECT 74.759 62.803 74.825 65.108 ;
      RECT 74.805 62.757 74.871 65.062 ;
      RECT 74.851 62.711 74.917 65.016 ;
      RECT 74.897 62.665 74.963 64.97 ;
      RECT 74.943 62.619 75.009 64.924 ;
      RECT 74.989 62.573 75.055 64.878 ;
      RECT 75.035 62.527 75.101 64.832 ;
      RECT 75.081 62.481 75.147 64.786 ;
      RECT 75.127 62.435 75.193 64.74 ;
      RECT 75.173 62.389 75.239 64.694 ;
      RECT 75.219 62.343 75.285 64.648 ;
      RECT 75.265 62.297 75.331 64.602 ;
      RECT 75.311 62.251 75.377 64.556 ;
      RECT 75.357 62.205 75.423 64.51 ;
      RECT 75.403 62.159 75.469 64.464 ;
      RECT 75.449 62.113 75.515 64.418 ;
      RECT 75.495 62.067 75.561 64.372 ;
      RECT 75.541 62.021 75.607 64.326 ;
      RECT 75.587 61.975 75.653 64.28 ;
      RECT 75.633 61.929 75.699 64.234 ;
      RECT 75.679 61.883 75.745 64.188 ;
      RECT 75.725 61.837 75.791 64.142 ;
      RECT 75.771 61.791 75.837 64.096 ;
      RECT 75.817 61.745 75.883 64.05 ;
      RECT 75.863 61.699 75.929 64.004 ;
      RECT 75.909 61.653 75.975 63.958 ;
      RECT 75.955 61.607 76.021 63.912 ;
      RECT 76.001 61.561 76.067 63.866 ;
      RECT 76.047 61.515 76.113 63.82 ;
      RECT 76.093 61.469 76.159 63.774 ;
      RECT 76.139 61.423 76.205 63.728 ;
      RECT 76.185 61.377 76.251 63.682 ;
      RECT 76.231 61.331 76.297 63.636 ;
      RECT 76.277 61.285 76.343 63.59 ;
      RECT 76.323 61.239 76.389 63.544 ;
      RECT 76.369 61.193 76.435 63.498 ;
      RECT 76.415 61.158 76.481 63.452 ;
      RECT 76.44 61.122 76.527 63.406 ;
      RECT 76.486 61.076 76.573 63.36 ;
      RECT 76.532 61.03 76.619 63.314 ;
      RECT 76.578 60.984 76.665 63.268 ;
      RECT 76.624 60.938 76.711 63.222 ;
      RECT 76.67 60.892 76.757 63.176 ;
      RECT 76.716 60.846 76.803 63.13 ;
      RECT 76.762 60.8 76.849 63.084 ;
      RECT 76.808 60.754 76.895 63.038 ;
      RECT 76.854 60.708 76.941 62.992 ;
      RECT 76.9 60.662 76.987 62.946 ;
      RECT 76.946 60.616 77.033 62.9 ;
      RECT 76.992 60.57 77.079 62.854 ;
      RECT 77.038 60.524 77.125 62.808 ;
      RECT 77.084 60.478 77.171 62.762 ;
      RECT 77.13 60.432 77.217 62.716 ;
      RECT 77.176 60.386 77.263 62.67 ;
      RECT 77.222 60.34 77.309 62.624 ;
      RECT 77.268 60.294 77.355 62.578 ;
      RECT 77.314 60.248 77.401 62.532 ;
      RECT 77.36 60.202 77.447 62.486 ;
      RECT 77.406 60.156 77.493 62.44 ;
      RECT 77.452 60.11 77.539 62.394 ;
      RECT 77.498 60.064 77.585 62.348 ;
      RECT 77.544 60.018 77.631 62.302 ;
      RECT 77.59 59.972 77.677 62.256 ;
      RECT 77.636 59.926 77.723 62.21 ;
      RECT 77.682 59.88 77.769 62.164 ;
      RECT 77.728 59.834 77.815 62.118 ;
      RECT 77.774 59.788 77.861 62.072 ;
      RECT 77.82 59.742 77.907 62.026 ;
      RECT 77.866 59.696 77.953 61.98 ;
      RECT 77.912 59.65 77.999 61.934 ;
      RECT 77.958 59.604 78.045 61.888 ;
      RECT 78.004 59.558 78.091 61.842 ;
      RECT 78.05 59.512 78.137 61.796 ;
      RECT 78.096 59.466 78.183 61.75 ;
      RECT 78.142 59.42 78.229 61.704 ;
      RECT 78.188 59.374 78.275 61.658 ;
      RECT 78.234 59.328 78.321 61.612 ;
      RECT 78.28 59.282 78.367 61.566 ;
      RECT 78.326 59.236 78.413 61.52 ;
      RECT 78.372 59.19 78.459 61.474 ;
      RECT 78.418 59.144 78.505 61.428 ;
      RECT 78.464 59.098 78.551 61.382 ;
      RECT 78.51 59.052 78.597 61.336 ;
      RECT 78.556 59.006 78.643 61.29 ;
      RECT 78.602 58.96 78.689 61.244 ;
      RECT 78.648 58.914 78.735 61.198 ;
      RECT 78.694 58.868 78.781 61.152 ;
      RECT 78.74 58.822 78.827 61.106 ;
      RECT 78.786 58.776 78.873 61.06 ;
      RECT 78.832 58.73 78.919 61.014 ;
      RECT 78.878 58.684 78.965 60.968 ;
      RECT 78.924 58.638 79.011 60.922 ;
      RECT 78.97 58.592 79.057 60.876 ;
      RECT 79.016 58.546 79.103 60.83 ;
      RECT 79.062 58.5 79.149 60.784 ;
      RECT 79.108 58.454 79.195 60.738 ;
      RECT 79.154 58.408 79.241 60.692 ;
      RECT 79.2 58.362 79.287 60.646 ;
      RECT 79.246 58.316 79.333 60.6 ;
      RECT 79.292 58.27 79.379 60.554 ;
      RECT 79.338 58.224 79.425 60.508 ;
      RECT 79.384 58.178 79.471 60.462 ;
      RECT 79.43 58.132 79.517 60.416 ;
      RECT 79.476 58.086 79.563 60.37 ;
      RECT 79.522 58.04 79.609 60.324 ;
      RECT 79.568 57.994 79.655 60.278 ;
      RECT 79.614 57.948 79.701 60.232 ;
      RECT 79.66 57.902 79.747 60.186 ;
      RECT 79.706 57.856 79.793 60.14 ;
      RECT 79.752 57.81 79.839 60.094 ;
      RECT 79.798 57.764 79.885 60.048 ;
      RECT 79.844 57.718 79.931 60.002 ;
      RECT 79.89 57.672 79.977 59.956 ;
      RECT 79.936 57.626 80.023 59.91 ;
      RECT 79.982 57.58 80.069 59.864 ;
      RECT 80.028 57.534 80.115 59.818 ;
      RECT 80.074 57.488 80.161 59.772 ;
      RECT 80.12 57.442 80.207 59.726 ;
      RECT 80.166 57.396 80.253 59.68 ;
      RECT 80.212 57.35 80.299 59.634 ;
      RECT 80.258 57.304 80.345 59.588 ;
      RECT 80.304 57.258 80.391 59.542 ;
      RECT 80.35 57.212 80.437 59.496 ;
      RECT 80.396 57.166 80.483 59.45 ;
      RECT 80.442 57.12 80.529 59.404 ;
      RECT 80.488 57.074 80.575 59.358 ;
      RECT 80.534 57.028 80.621 59.312 ;
      RECT 80.58 56.982 80.667 59.266 ;
      RECT 80.626 56.936 80.713 59.22 ;
      RECT 80.672 56.89 80.759 59.174 ;
      RECT 80.718 56.844 80.805 59.128 ;
      RECT 80.764 56.798 80.851 59.082 ;
      RECT 80.81 56.752 80.897 59.036 ;
      RECT 80.856 56.706 80.943 58.99 ;
      RECT 80.902 56.66 80.989 58.944 ;
      RECT 80.948 56.614 81.035 58.898 ;
      RECT 80.994 56.568 81.081 58.852 ;
      RECT 81.04 56.522 81.127 58.806 ;
      RECT 81.086 56.476 81.173 58.76 ;
      RECT 81.132 56.43 81.219 58.714 ;
      RECT 81.178 56.384 81.265 58.668 ;
      RECT 81.224 56.338 81.311 58.622 ;
      RECT 81.27 56.292 81.357 58.576 ;
      RECT 81.316 56.246 81.403 58.53 ;
      RECT 81.362 56.199 81.449 58.484 ;
      RECT 81.408 56.175 81.495 58.438 ;
      RECT 81.408 56.175 81.541 58.392 ;
      RECT 81.408 56.175 81.587 58.346 ;
      RECT 81.408 56.175 81.633 58.3 ;
      RECT 81.408 56.175 81.679 58.254 ;
      RECT 81.408 56.175 81.725 58.208 ;
      RECT 81.408 56.175 81.771 58.162 ;
      RECT 81.408 56.175 81.817 58.116 ;
      RECT 81.408 56.175 81.863 58.07 ;
      RECT 81.408 56.175 81.909 58.024 ;
      RECT 81.408 56.175 81.955 57.978 ;
      RECT 81.408 56.175 82.001 57.932 ;
      RECT 81.408 56.175 82.047 57.886 ;
      RECT 81.408 56.175 82.093 57.84 ;
      RECT 81.408 56.175 82.139 57.794 ;
      RECT 81.408 56.175 82.185 57.748 ;
      RECT 81.408 56.175 82.231 57.702 ;
      RECT 81.408 56.175 82.277 57.656 ;
      RECT 81.408 56.175 82.323 57.61 ;
      RECT 81.408 56.175 82.369 57.564 ;
      RECT 81.408 56.175 82.415 57.518 ;
      RECT 81.408 56.175 82.461 57.472 ;
      RECT 81.408 56.175 82.507 57.426 ;
      RECT 81.408 56.175 82.553 57.38 ;
      RECT 80.258 57.304 82.585 57.341 ;
      RECT 81.408 56.175 110 57.325 ;
      RECT 63.675 85.392 68.325 110 ;
      RECT 63.675 85.392 68.371 88.167 ;
      RECT 63.675 85.392 68.417 88.121 ;
      RECT 63.675 85.392 68.463 88.075 ;
      RECT 63.675 85.392 68.509 88.029 ;
      RECT 63.675 85.392 68.555 87.983 ;
      RECT 63.675 85.392 68.601 87.937 ;
      RECT 63.675 85.392 68.647 87.891 ;
      RECT 63.675 85.392 68.693 87.845 ;
      RECT 63.675 85.392 68.739 87.799 ;
      RECT 63.675 85.392 68.785 87.753 ;
      RECT 63.675 85.392 68.831 87.707 ;
      RECT 63.675 85.392 68.877 87.661 ;
      RECT 63.675 85.392 68.923 87.615 ;
      RECT 63.675 85.392 68.969 87.569 ;
      RECT 63.675 85.392 69.015 87.523 ;
      RECT 63.675 85.392 69.061 87.477 ;
      RECT 63.675 85.392 69.107 87.431 ;
      RECT 63.675 85.392 69.153 87.385 ;
      RECT 63.675 85.392 69.199 87.339 ;
      RECT 63.675 85.392 69.245 87.293 ;
      RECT 63.675 85.392 69.291 87.247 ;
      RECT 63.675 85.392 69.337 87.201 ;
      RECT 63.675 85.392 69.383 87.155 ;
      RECT 63.675 85.392 69.429 87.109 ;
      RECT 63.675 85.392 69.475 87.063 ;
      RECT 63.675 85.392 69.521 87.017 ;
      RECT 63.675 85.392 69.567 86.971 ;
      RECT 63.675 85.392 69.613 86.925 ;
      RECT 63.675 85.392 69.659 86.879 ;
      RECT 63.675 85.392 69.705 86.833 ;
      RECT 63.675 85.392 69.751 86.787 ;
      RECT 63.675 85.392 69.797 86.741 ;
      RECT 63.675 85.392 69.843 86.695 ;
      RECT 63.675 85.392 69.889 86.649 ;
      RECT 63.675 85.392 69.935 86.603 ;
      RECT 63.675 85.392 69.981 86.557 ;
      RECT 63.675 85.392 70.027 86.511 ;
      RECT 63.675 85.392 70.073 86.465 ;
      RECT 63.675 85.392 70.119 86.419 ;
      RECT 63.675 85.392 70.165 86.373 ;
      RECT 63.675 85.392 70.211 86.327 ;
      RECT 63.675 85.392 70.257 86.281 ;
      RECT 63.675 85.392 70.303 86.235 ;
      RECT 63.675 85.392 70.349 86.189 ;
      RECT 63.675 85.392 70.395 86.143 ;
      RECT 63.675 85.392 70.441 86.097 ;
      RECT 63.675 85.392 70.487 86.051 ;
      RECT 63.675 85.392 70.533 86.005 ;
      RECT 63.675 85.392 70.579 85.959 ;
      RECT 63.675 85.392 70.625 85.913 ;
      RECT 63.675 85.392 70.671 85.867 ;
      RECT 63.675 85.392 70.717 85.821 ;
      RECT 63.675 85.392 70.763 85.775 ;
      RECT 63.675 85.392 70.809 85.729 ;
      RECT 63.675 85.392 70.855 85.683 ;
      RECT 63.675 85.392 70.901 85.637 ;
      RECT 63.675 85.392 70.947 85.591 ;
      RECT 63.675 85.392 70.993 85.545 ;
      RECT 63.675 85.392 71.039 85.499 ;
      RECT 63.721 85.346 71.131 85.407 ;
      RECT 71.081 77.986 71.131 85.407 ;
      RECT 63.767 85.3 71.177 85.361 ;
      RECT 71.127 77.94 71.177 85.361 ;
      RECT 63.813 85.254 71.223 85.315 ;
      RECT 71.173 77.894 71.223 85.315 ;
      RECT 63.859 85.208 71.269 85.269 ;
      RECT 71.219 77.848 71.269 85.269 ;
      RECT 63.905 85.162 71.315 85.223 ;
      RECT 71.265 77.802 71.315 85.223 ;
      RECT 63.951 85.116 71.361 85.177 ;
      RECT 71.311 77.756 71.361 85.177 ;
      RECT 63.997 85.07 71.407 85.131 ;
      RECT 71.357 77.71 71.407 85.131 ;
      RECT 64.043 85.024 71.453 85.085 ;
      RECT 71.403 77.664 71.453 85.085 ;
      RECT 64.089 84.978 71.499 85.039 ;
      RECT 71.449 77.618 71.499 85.039 ;
      RECT 64.135 84.932 71.545 84.993 ;
      RECT 71.495 77.572 71.545 84.993 ;
      RECT 64.181 84.886 71.591 84.947 ;
      RECT 71.541 77.526 71.591 84.947 ;
      RECT 64.227 84.84 71.637 84.901 ;
      RECT 71.587 77.48 71.637 84.901 ;
      RECT 64.273 84.794 71.683 84.855 ;
      RECT 71.633 77.434 71.683 84.855 ;
      RECT 64.319 84.748 71.729 84.809 ;
      RECT 71.679 77.388 71.729 84.809 ;
      RECT 64.365 84.702 71.775 84.763 ;
      RECT 71.725 77.342 71.775 84.763 ;
      RECT 64.411 84.656 71.821 84.717 ;
      RECT 71.771 77.296 71.821 84.717 ;
      RECT 64.457 84.61 71.867 84.671 ;
      RECT 71.817 77.25 71.867 84.671 ;
      RECT 64.503 84.564 71.913 84.625 ;
      RECT 71.863 77.204 71.913 84.625 ;
      RECT 64.549 84.518 71.959 84.579 ;
      RECT 71.909 77.158 71.959 84.579 ;
      RECT 64.595 84.472 72.005 84.533 ;
      RECT 71.955 77.112 72.005 84.533 ;
      RECT 64.641 84.426 72.051 84.487 ;
      RECT 72.001 77.066 72.051 84.487 ;
      RECT 64.687 84.38 72.097 84.441 ;
      RECT 72.047 77.02 72.097 84.441 ;
      RECT 64.733 84.334 72.143 84.395 ;
      RECT 72.093 76.974 72.143 84.395 ;
      RECT 64.779 84.288 72.189 84.349 ;
      RECT 72.139 76.928 72.189 84.349 ;
      RECT 64.825 84.242 72.235 84.303 ;
      RECT 72.185 76.882 72.235 84.303 ;
      RECT 64.871 84.196 72.281 84.257 ;
      RECT 72.231 76.836 72.281 84.257 ;
      RECT 64.917 84.15 72.327 84.211 ;
      RECT 72.277 76.79 72.327 84.211 ;
      RECT 64.963 84.104 72.373 84.165 ;
      RECT 72.323 76.744 72.373 84.165 ;
      RECT 65.009 84.058 72.419 84.119 ;
      RECT 72.369 76.698 72.419 84.119 ;
      RECT 65.055 84.012 72.465 84.073 ;
      RECT 72.415 76.652 72.465 84.073 ;
      RECT 65.101 83.966 72.511 84.027 ;
      RECT 72.461 76.606 72.511 84.027 ;
      RECT 65.147 83.92 72.557 83.981 ;
      RECT 72.507 76.56 72.557 83.981 ;
      RECT 65.193 83.874 72.603 83.935 ;
      RECT 72.553 76.514 72.603 83.935 ;
      RECT 65.239 83.828 72.649 83.889 ;
      RECT 72.599 76.468 72.649 83.889 ;
      RECT 65.285 83.782 72.695 83.843 ;
      RECT 72.645 76.422 72.695 83.843 ;
      RECT 65.331 83.736 72.741 83.797 ;
      RECT 72.691 76.376 72.741 83.797 ;
      RECT 65.377 83.69 72.787 83.751 ;
      RECT 72.737 76.33 72.787 83.751 ;
      RECT 65.423 83.644 72.833 83.705 ;
      RECT 72.783 76.284 72.833 83.705 ;
      RECT 65.469 83.598 72.879 83.659 ;
      RECT 72.829 76.238 72.879 83.659 ;
      RECT 65.515 83.552 72.925 83.613 ;
      RECT 72.875 76.192 72.925 83.613 ;
      RECT 65.561 83.506 72.971 83.567 ;
      RECT 72.921 76.146 72.971 83.567 ;
      RECT 65.607 83.46 73.017 83.521 ;
      RECT 72.967 76.1 73.017 83.521 ;
      RECT 65.653 83.414 73.063 83.475 ;
      RECT 73.013 76.054 73.063 83.475 ;
      RECT 65.699 83.368 73.109 83.429 ;
      RECT 73.059 76.008 73.109 83.429 ;
      RECT 65.745 83.322 73.155 83.383 ;
      RECT 73.105 75.962 73.155 83.383 ;
      RECT 65.791 83.276 73.201 83.337 ;
      RECT 73.151 75.916 73.201 83.337 ;
      RECT 65.837 83.23 73.247 83.291 ;
      RECT 73.197 75.87 73.247 83.291 ;
      RECT 65.883 83.184 73.293 83.245 ;
      RECT 73.243 75.824 73.293 83.245 ;
      RECT 65.929 83.138 73.339 83.199 ;
      RECT 73.289 75.778 73.339 83.199 ;
      RECT 65.975 83.092 73.385 83.153 ;
      RECT 73.335 75.732 73.385 83.153 ;
      RECT 66.021 83.046 73.431 83.107 ;
      RECT 73.381 75.686 73.431 83.107 ;
      RECT 66.067 83 73.477 83.061 ;
      RECT 73.427 75.64 73.477 83.061 ;
      RECT 66.113 82.954 73.523 83.015 ;
      RECT 73.473 75.594 73.523 83.015 ;
      RECT 66.159 82.908 73.569 82.969 ;
      RECT 73.519 75.548 73.569 82.969 ;
      RECT 66.205 82.862 73.615 82.923 ;
      RECT 73.565 75.502 73.615 82.923 ;
      RECT 66.251 82.816 73.661 82.877 ;
      RECT 73.611 75.456 73.661 82.877 ;
      RECT 66.297 82.77 73.707 82.831 ;
      RECT 73.657 75.41 73.707 82.831 ;
      RECT 66.343 82.724 73.753 82.785 ;
      RECT 73.703 75.364 73.753 82.785 ;
      RECT 66.389 82.678 73.799 82.739 ;
      RECT 73.749 75.318 73.799 82.739 ;
      RECT 66.435 82.632 73.845 82.693 ;
      RECT 73.795 75.272 73.845 82.693 ;
      RECT 66.481 82.586 73.891 82.647 ;
      RECT 73.841 75.226 73.891 82.647 ;
      RECT 66.527 82.54 73.937 82.601 ;
      RECT 73.887 75.18 73.937 82.601 ;
      RECT 66.573 82.494 73.983 82.555 ;
      RECT 73.933 75.134 73.983 82.555 ;
      RECT 66.619 82.448 74.029 82.509 ;
      RECT 73.979 75.088 74.029 82.509 ;
      RECT 66.665 82.402 74.075 82.463 ;
      RECT 74.025 75.042 74.075 82.463 ;
      RECT 66.711 82.356 74.121 82.417 ;
      RECT 74.071 74.996 74.121 82.417 ;
      RECT 66.757 82.31 74.167 82.371 ;
      RECT 74.117 74.95 74.167 82.371 ;
      RECT 66.803 82.264 74.213 82.325 ;
      RECT 74.163 74.904 74.213 82.325 ;
      RECT 66.849 82.218 74.259 82.279 ;
      RECT 74.209 74.858 74.259 82.279 ;
      RECT 66.895 82.172 74.305 82.233 ;
      RECT 74.255 74.812 74.305 82.233 ;
      RECT 66.941 82.126 74.351 82.187 ;
      RECT 74.301 74.766 74.351 82.187 ;
      RECT 66.987 82.08 74.397 82.141 ;
      RECT 74.347 74.72 74.397 82.141 ;
      RECT 67.033 82.034 74.443 82.095 ;
      RECT 74.393 74.674 74.443 82.095 ;
      RECT 67.079 81.988 74.489 82.049 ;
      RECT 74.439 74.628 74.489 82.049 ;
      RECT 67.125 81.942 74.535 82.003 ;
      RECT 74.485 74.582 74.535 82.003 ;
      RECT 67.171 81.896 74.581 81.957 ;
      RECT 74.531 74.536 74.581 81.957 ;
      RECT 67.217 81.85 74.627 81.911 ;
      RECT 74.577 74.49 74.627 81.911 ;
      RECT 67.263 81.804 74.673 81.865 ;
      RECT 74.623 74.444 74.673 81.865 ;
      RECT 67.309 81.758 74.719 81.819 ;
      RECT 74.669 74.398 74.719 81.819 ;
      RECT 67.355 81.712 74.765 81.773 ;
      RECT 74.715 74.352 74.765 81.773 ;
      RECT 67.401 81.666 74.811 81.727 ;
      RECT 74.761 74.306 74.811 81.727 ;
      RECT 67.447 81.62 74.857 81.681 ;
      RECT 74.807 74.26 74.857 81.681 ;
      RECT 67.493 81.574 74.903 81.635 ;
      RECT 74.853 74.214 74.903 81.635 ;
      RECT 67.539 81.528 74.949 81.589 ;
      RECT 74.899 74.168 74.949 81.589 ;
      RECT 67.585 81.482 74.995 81.543 ;
      RECT 74.945 74.122 74.995 81.543 ;
      RECT 67.631 81.436 75.041 81.497 ;
      RECT 74.991 74.076 75.041 81.497 ;
      RECT 67.677 81.39 75.087 81.451 ;
      RECT 75.037 74.03 75.087 81.451 ;
      RECT 67.723 81.344 75.133 81.405 ;
      RECT 75.083 73.984 75.133 81.405 ;
      RECT 67.769 81.298 75.179 81.359 ;
      RECT 75.129 73.938 75.179 81.359 ;
      RECT 67.815 81.252 75.225 81.313 ;
      RECT 75.175 73.892 75.225 81.313 ;
      RECT 67.861 81.206 75.271 81.267 ;
      RECT 75.221 73.846 75.271 81.267 ;
      RECT 67.907 81.16 75.317 81.221 ;
      RECT 75.267 73.8 75.317 81.221 ;
      RECT 67.953 81.114 75.363 81.175 ;
      RECT 75.313 73.754 75.363 81.175 ;
      RECT 67.999 81.068 75.409 81.129 ;
      RECT 75.359 73.708 75.409 81.129 ;
      RECT 68.045 81.022 75.455 81.083 ;
      RECT 75.405 73.662 75.455 81.083 ;
      RECT 68.091 80.976 75.501 81.037 ;
      RECT 75.451 73.616 75.501 81.037 ;
      RECT 68.137 80.93 75.547 80.991 ;
      RECT 75.497 73.57 75.547 80.991 ;
      RECT 68.183 80.884 75.593 80.945 ;
      RECT 75.543 73.524 75.593 80.945 ;
      RECT 68.229 80.838 75.639 80.899 ;
      RECT 75.589 73.478 75.639 80.899 ;
      RECT 68.275 80.792 75.685 80.853 ;
      RECT 75.635 73.432 75.685 80.853 ;
      RECT 68.321 80.746 75.731 80.807 ;
      RECT 75.681 73.386 75.731 80.807 ;
      RECT 68.367 80.7 75.777 80.761 ;
      RECT 75.727 73.34 75.777 80.761 ;
      RECT 68.413 80.654 75.823 80.715 ;
      RECT 75.773 73.294 75.823 80.715 ;
      RECT 68.459 80.608 75.869 80.669 ;
      RECT 75.819 73.248 75.869 80.669 ;
      RECT 68.505 80.562 75.915 80.623 ;
      RECT 75.865 73.202 75.915 80.623 ;
      RECT 68.551 80.516 75.961 80.577 ;
      RECT 75.911 73.156 75.961 80.577 ;
      RECT 68.597 80.47 76.007 80.531 ;
      RECT 75.957 73.11 76.007 80.531 ;
      RECT 68.643 80.424 76.053 80.485 ;
      RECT 76.003 73.064 76.053 80.485 ;
      RECT 68.689 80.378 76.099 80.439 ;
      RECT 76.049 73.018 76.099 80.439 ;
      RECT 68.735 80.332 76.145 80.393 ;
      RECT 76.095 72.972 76.145 80.393 ;
      RECT 68.781 80.286 76.191 80.347 ;
      RECT 76.141 72.926 76.191 80.347 ;
      RECT 68.827 80.24 76.237 80.301 ;
      RECT 76.187 72.88 76.237 80.301 ;
      RECT 68.873 80.194 76.283 80.255 ;
      RECT 76.233 72.834 76.283 80.255 ;
      RECT 68.919 80.148 76.329 80.209 ;
      RECT 76.279 72.788 76.329 80.209 ;
      RECT 68.965 80.102 76.375 80.163 ;
      RECT 76.325 72.742 76.375 80.163 ;
      RECT 69.011 80.056 76.421 80.117 ;
      RECT 76.371 72.696 76.421 80.117 ;
      RECT 69.057 80.01 76.467 80.071 ;
      RECT 76.417 72.65 76.467 80.071 ;
      RECT 69.103 79.964 76.513 80.025 ;
      RECT 76.463 72.604 76.513 80.025 ;
      RECT 69.149 79.918 76.559 79.979 ;
      RECT 76.509 72.558 76.559 79.979 ;
      RECT 69.195 79.872 76.605 79.933 ;
      RECT 76.555 72.512 76.605 79.933 ;
      RECT 69.241 79.826 76.651 79.887 ;
      RECT 76.601 72.466 76.651 79.887 ;
      RECT 69.287 79.78 76.697 79.841 ;
      RECT 76.647 72.42 76.697 79.841 ;
      RECT 69.333 79.734 76.743 79.795 ;
      RECT 76.693 72.374 76.743 79.795 ;
      RECT 69.379 79.688 76.789 79.749 ;
      RECT 76.739 72.328 76.789 79.749 ;
      RECT 69.425 79.642 76.825 79.708 ;
      RECT 71.035 78.032 71.085 85.453 ;
      RECT 69.471 79.596 76.871 79.667 ;
      RECT 76.785 72.282 76.871 79.667 ;
      RECT 69.517 79.55 76.917 79.621 ;
      RECT 76.831 72.236 76.917 79.621 ;
      RECT 69.563 79.504 76.963 79.575 ;
      RECT 76.877 72.19 76.963 79.575 ;
      RECT 69.609 79.458 77.009 79.529 ;
      RECT 76.923 72.144 77.009 79.529 ;
      RECT 69.655 79.412 77.055 79.483 ;
      RECT 76.969 72.098 77.055 79.483 ;
      RECT 69.701 79.366 77.101 79.437 ;
      RECT 77.015 72.052 77.101 79.437 ;
      RECT 69.747 79.32 77.147 79.391 ;
      RECT 77.061 72.006 77.147 79.391 ;
      RECT 69.793 79.274 77.193 79.345 ;
      RECT 77.107 71.96 77.193 79.345 ;
      RECT 69.839 79.228 77.239 79.299 ;
      RECT 77.153 71.914 77.239 79.299 ;
      RECT 69.885 79.182 77.285 79.253 ;
      RECT 77.199 71.868 77.285 79.253 ;
      RECT 69.931 79.136 77.331 79.207 ;
      RECT 77.245 71.822 77.331 79.207 ;
      RECT 69.977 79.09 77.377 79.161 ;
      RECT 77.291 71.776 77.377 79.161 ;
      RECT 70.023 79.044 77.423 79.115 ;
      RECT 77.337 71.73 77.423 79.115 ;
      RECT 70.069 78.998 77.469 79.069 ;
      RECT 77.383 71.684 77.469 79.069 ;
      RECT 70.115 78.952 77.515 79.023 ;
      RECT 77.429 71.638 77.515 79.023 ;
      RECT 70.161 78.906 77.561 78.977 ;
      RECT 77.475 71.592 77.561 78.977 ;
      RECT 70.207 78.86 77.607 78.931 ;
      RECT 77.521 71.546 77.607 78.931 ;
      RECT 70.253 78.814 77.653 78.885 ;
      RECT 77.567 71.5 77.653 78.885 ;
      RECT 70.299 78.768 77.699 78.839 ;
      RECT 77.613 71.454 77.699 78.839 ;
      RECT 70.345 78.722 77.745 78.793 ;
      RECT 77.659 71.408 77.745 78.793 ;
      RECT 70.391 78.676 77.791 78.747 ;
      RECT 77.705 71.362 77.791 78.747 ;
      RECT 70.437 78.63 77.837 78.701 ;
      RECT 77.751 71.316 77.837 78.701 ;
      RECT 70.483 78.584 77.883 78.655 ;
      RECT 77.797 71.27 77.883 78.655 ;
      RECT 70.529 78.538 77.929 78.609 ;
      RECT 77.843 71.224 77.929 78.609 ;
      RECT 70.575 78.492 77.975 78.563 ;
      RECT 77.889 71.178 77.975 78.563 ;
      RECT 70.621 78.446 78.021 78.517 ;
      RECT 77.935 71.132 78.021 78.517 ;
      RECT 70.667 78.4 78.067 78.471 ;
      RECT 77.981 71.086 78.067 78.471 ;
      RECT 70.713 78.354 78.113 78.425 ;
      RECT 78.027 71.04 78.113 78.425 ;
      RECT 70.759 78.308 78.159 78.379 ;
      RECT 78.073 70.994 78.159 78.379 ;
      RECT 70.805 78.262 78.205 78.333 ;
      RECT 78.119 70.948 78.205 78.333 ;
      RECT 70.851 78.216 78.251 78.287 ;
      RECT 78.165 70.902 78.251 78.287 ;
      RECT 70.897 78.17 78.297 78.241 ;
      RECT 78.211 70.856 78.297 78.241 ;
      RECT 70.943 78.124 78.343 78.195 ;
      RECT 78.257 70.81 78.343 78.195 ;
      RECT 70.989 78.078 78.389 78.149 ;
      RECT 78.303 70.764 78.389 78.149 ;
      RECT 78.349 70.718 78.435 78.103 ;
      RECT 78.395 70.672 78.481 78.057 ;
      RECT 78.441 70.626 78.527 78.011 ;
      RECT 78.487 70.58 78.573 77.965 ;
      RECT 78.533 70.534 78.619 77.919 ;
      RECT 78.579 70.488 78.665 77.873 ;
      RECT 78.625 70.442 78.711 77.827 ;
      RECT 78.671 70.396 78.757 77.781 ;
      RECT 78.717 70.35 78.803 77.735 ;
      RECT 78.763 70.304 78.849 77.689 ;
      RECT 78.809 70.258 78.895 77.643 ;
      RECT 78.855 70.212 78.941 77.597 ;
      RECT 78.901 70.166 78.987 77.551 ;
      RECT 78.947 70.12 79.033 77.505 ;
      RECT 78.993 70.074 79.079 77.459 ;
      RECT 79.039 70.028 79.125 77.413 ;
      RECT 79.085 69.982 79.171 77.367 ;
      RECT 79.131 69.936 79.217 77.321 ;
      RECT 79.177 69.89 79.263 77.275 ;
      RECT 79.223 69.844 79.309 77.229 ;
      RECT 79.269 69.798 79.355 77.183 ;
      RECT 79.315 69.752 79.401 77.137 ;
      RECT 79.361 69.706 79.447 77.091 ;
      RECT 79.407 69.66 79.493 77.045 ;
      RECT 79.453 69.614 79.539 76.999 ;
      RECT 79.499 69.568 79.585 76.953 ;
      RECT 79.545 69.522 79.631 76.907 ;
      RECT 79.591 69.476 79.677 76.861 ;
      RECT 79.637 69.43 79.723 76.815 ;
      RECT 79.683 69.384 79.769 76.769 ;
      RECT 79.729 69.338 79.815 76.723 ;
      RECT 79.775 69.292 79.861 76.677 ;
      RECT 79.821 69.246 79.907 76.631 ;
      RECT 79.867 69.2 79.953 76.585 ;
      RECT 79.913 69.154 79.999 76.539 ;
      RECT 79.959 69.108 80.045 76.493 ;
      RECT 80.005 69.062 80.091 76.447 ;
      RECT 80.051 69.016 80.137 76.401 ;
      RECT 80.097 68.97 80.183 76.355 ;
      RECT 80.143 68.924 80.229 76.309 ;
      RECT 80.189 68.878 80.275 76.263 ;
      RECT 80.235 68.832 80.321 76.217 ;
      RECT 80.281 68.786 80.367 76.171 ;
      RECT 80.327 68.74 80.413 76.125 ;
      RECT 80.373 68.694 80.459 76.079 ;
      RECT 80.419 68.648 80.505 76.033 ;
      RECT 80.465 68.602 80.551 75.987 ;
      RECT 80.511 68.556 80.597 75.941 ;
      RECT 80.557 68.51 80.643 75.895 ;
      RECT 80.603 68.464 80.689 75.849 ;
      RECT 80.649 68.418 80.735 75.803 ;
      RECT 80.695 68.372 80.781 75.757 ;
      RECT 80.741 68.326 80.827 75.711 ;
      RECT 80.787 68.28 80.873 75.665 ;
      RECT 80.833 68.234 80.919 75.619 ;
      RECT 80.879 68.188 80.965 75.573 ;
      RECT 80.925 68.142 81.011 75.527 ;
      RECT 80.971 68.096 81.057 75.481 ;
      RECT 81.017 68.05 81.103 75.435 ;
      RECT 81.063 68.004 81.149 75.389 ;
      RECT 81.109 67.958 81.195 75.343 ;
      RECT 81.155 67.912 81.241 75.297 ;
      RECT 81.201 67.866 81.287 75.251 ;
      RECT 81.247 67.82 81.333 75.205 ;
      RECT 81.293 67.774 81.379 75.159 ;
      RECT 81.339 67.728 81.425 75.113 ;
      RECT 81.385 67.682 81.471 75.067 ;
      RECT 81.431 67.636 81.517 75.021 ;
      RECT 81.477 67.59 81.563 74.975 ;
      RECT 81.523 67.544 81.609 74.929 ;
      RECT 81.569 67.498 81.655 74.883 ;
      RECT 81.615 67.452 81.701 74.837 ;
      RECT 81.661 67.406 81.747 74.791 ;
      RECT 81.707 67.36 81.793 74.745 ;
      RECT 81.753 67.314 81.839 74.699 ;
      RECT 81.799 67.268 81.885 74.653 ;
      RECT 81.845 67.222 81.931 74.607 ;
      RECT 81.891 67.176 81.977 74.561 ;
      RECT 81.937 67.13 82.023 74.515 ;
      RECT 81.983 67.084 82.069 74.469 ;
      RECT 82.029 67.038 82.115 74.423 ;
      RECT 82.075 66.992 82.161 74.377 ;
      RECT 82.121 66.946 82.207 74.331 ;
      RECT 82.167 66.9 82.253 74.285 ;
      RECT 82.213 66.854 82.299 74.239 ;
      RECT 82.259 66.808 82.345 74.193 ;
      RECT 82.305 66.762 82.391 74.147 ;
      RECT 82.351 66.716 82.437 74.101 ;
      RECT 82.397 66.67 82.483 74.055 ;
      RECT 82.443 66.624 82.529 74.009 ;
      RECT 82.489 66.578 82.575 73.963 ;
      RECT 82.535 66.532 82.621 73.917 ;
      RECT 82.581 66.486 82.667 73.871 ;
      RECT 82.627 66.44 82.713 73.825 ;
      RECT 82.673 66.394 82.759 73.779 ;
      RECT 82.719 66.348 82.805 73.733 ;
      RECT 82.765 66.302 82.851 73.687 ;
      RECT 82.811 66.256 82.897 73.641 ;
      RECT 82.903 66.171 82.943 73.595 ;
      RECT 82.935 66.132 82.989 73.549 ;
      RECT 82.981 66.086 83.035 73.503 ;
      RECT 83.027 66.04 83.081 73.457 ;
      RECT 83.073 65.994 83.127 73.411 ;
      RECT 83.119 65.948 83.173 73.365 ;
      RECT 83.165 65.902 83.219 73.319 ;
      RECT 83.211 65.856 83.265 73.273 ;
      RECT 83.257 65.81 83.311 73.227 ;
      RECT 83.303 65.764 83.357 73.181 ;
      RECT 83.349 65.718 83.403 73.135 ;
      RECT 83.395 65.672 83.449 73.089 ;
      RECT 83.441 65.626 83.495 73.043 ;
      RECT 83.487 65.58 83.541 72.997 ;
      RECT 83.533 65.534 83.587 72.951 ;
      RECT 83.579 65.488 83.633 72.905 ;
      RECT 83.625 65.442 83.679 72.859 ;
      RECT 83.671 65.396 83.725 72.813 ;
      RECT 83.717 65.35 83.771 72.767 ;
      RECT 83.763 65.304 83.817 72.721 ;
      RECT 83.809 65.258 83.863 72.675 ;
      RECT 83.855 65.212 83.909 72.629 ;
      RECT 83.901 65.166 83.955 72.583 ;
      RECT 83.947 65.12 84.001 72.537 ;
      RECT 83.993 65.074 84.047 72.491 ;
      RECT 84.039 65.028 84.093 72.445 ;
      RECT 84.085 64.982 84.139 72.399 ;
      RECT 84.131 64.936 84.185 72.353 ;
      RECT 84.177 64.89 84.231 72.307 ;
      RECT 84.223 64.844 84.277 72.261 ;
      RECT 84.269 64.798 84.323 72.215 ;
      RECT 84.315 64.752 84.369 72.169 ;
      RECT 84.361 64.706 84.415 72.123 ;
      RECT 84.407 64.66 84.461 72.077 ;
      RECT 84.453 64.614 84.507 72.031 ;
      RECT 84.499 64.568 84.553 71.985 ;
      RECT 84.545 64.522 84.599 71.939 ;
      RECT 84.591 64.476 84.645 71.893 ;
      RECT 84.637 64.43 84.691 71.847 ;
      RECT 84.683 64.384 84.737 71.801 ;
      RECT 84.729 64.338 84.783 71.755 ;
      RECT 84.775 64.292 84.829 71.709 ;
      RECT 84.821 64.246 84.875 71.663 ;
      RECT 84.867 64.2 84.921 71.617 ;
      RECT 84.913 64.154 84.967 71.571 ;
      RECT 84.959 64.108 85.013 71.525 ;
      RECT 85.005 64.062 85.059 71.479 ;
      RECT 85.051 64.016 85.105 71.433 ;
      RECT 85.097 63.97 85.151 71.387 ;
      RECT 85.143 63.924 85.197 71.341 ;
      RECT 85.189 63.878 85.243 71.295 ;
      RECT 85.235 63.832 85.289 71.249 ;
      RECT 85.281 63.786 85.335 71.203 ;
      RECT 85.327 63.74 85.381 71.157 ;
      RECT 85.373 63.696 85.427 71.111 ;
      RECT 85.415 63.675 85.473 71.065 ;
      RECT 82.857 66.21 82.943 73.595 ;
      RECT 85.415 63.675 85.519 71.019 ;
      RECT 85.415 63.675 85.565 70.973 ;
      RECT 85.415 63.675 85.611 70.927 ;
      RECT 85.415 63.675 85.657 70.881 ;
      RECT 85.415 63.675 85.703 70.835 ;
      RECT 85.415 63.675 85.749 70.789 ;
      RECT 85.415 63.675 85.795 70.743 ;
      RECT 85.415 63.675 85.841 70.697 ;
      RECT 85.415 63.675 85.887 70.651 ;
      RECT 85.415 63.675 85.933 70.605 ;
      RECT 85.415 63.675 85.979 70.559 ;
      RECT 85.415 63.675 86.025 70.513 ;
      RECT 85.415 63.675 86.071 70.467 ;
      RECT 85.415 63.675 86.117 70.421 ;
      RECT 85.415 63.675 86.163 70.375 ;
      RECT 85.415 63.675 86.209 70.329 ;
      RECT 85.415 63.675 86.255 70.283 ;
      RECT 85.415 63.675 86.301 70.237 ;
      RECT 85.415 63.675 86.347 70.191 ;
      RECT 85.415 63.675 86.393 70.145 ;
      RECT 85.415 63.675 86.439 70.099 ;
      RECT 85.415 63.675 86.485 70.053 ;
      RECT 85.415 63.675 86.531 70.007 ;
      RECT 85.415 63.675 86.577 69.961 ;
      RECT 85.415 63.675 86.623 69.915 ;
      RECT 85.415 63.675 86.669 69.869 ;
      RECT 85.415 63.675 86.715 69.823 ;
      RECT 85.415 63.675 86.761 69.777 ;
      RECT 85.415 63.675 86.807 69.731 ;
      RECT 85.415 63.675 86.853 69.685 ;
      RECT 85.415 63.675 86.899 69.639 ;
      RECT 85.415 63.675 86.945 69.593 ;
      RECT 85.415 63.675 86.991 69.547 ;
      RECT 85.415 63.675 87.037 69.501 ;
      RECT 85.415 63.675 87.083 69.455 ;
      RECT 85.415 63.675 87.129 69.409 ;
      RECT 85.415 63.675 87.175 69.363 ;
      RECT 85.415 63.675 87.221 69.317 ;
      RECT 85.415 63.675 87.267 69.271 ;
      RECT 85.415 63.675 87.313 69.225 ;
      RECT 85.415 63.675 87.359 69.179 ;
      RECT 85.415 63.675 87.405 69.133 ;
      RECT 85.415 63.675 87.451 69.087 ;
      RECT 85.415 63.675 87.497 69.041 ;
      RECT 85.415 63.675 87.543 68.995 ;
      RECT 85.415 63.675 87.589 68.949 ;
      RECT 85.415 63.675 87.635 68.903 ;
      RECT 85.415 63.675 87.681 68.857 ;
      RECT 85.415 63.675 87.727 68.811 ;
      RECT 85.415 63.675 87.773 68.765 ;
      RECT 85.415 63.675 87.819 68.719 ;
      RECT 85.415 63.675 87.865 68.673 ;
      RECT 85.415 63.675 87.911 68.627 ;
      RECT 85.415 63.675 87.957 68.581 ;
      RECT 85.415 63.675 88.003 68.535 ;
      RECT 85.415 63.675 88.049 68.489 ;
      RECT 85.415 63.675 88.095 68.443 ;
      RECT 85.415 63.675 88.141 68.397 ;
      RECT 80.741 68.326 88.187 68.351 ;
      RECT 85.415 63.675 88.19 68.326 ;
      RECT 85.415 63.675 110 68.325 ;
      RECT 77.175 92.037 78.325 110 ;
      RECT 77.175 92.037 78.371 92.272 ;
      RECT 77.175 92.037 78.417 92.226 ;
      RECT 77.175 92.037 78.463 92.18 ;
      RECT 77.175 92.037 78.509 92.134 ;
      RECT 77.175 92.037 78.555 92.088 ;
      RECT 77.221 91.991 78.601 92.042 ;
      RECT 77.267 91.945 78.647 91.996 ;
      RECT 77.313 91.899 78.693 91.95 ;
      RECT 77.359 91.853 78.739 91.904 ;
      RECT 77.405 91.807 78.785 91.858 ;
      RECT 77.451 91.761 78.831 91.812 ;
      RECT 77.497 91.715 78.877 91.766 ;
      RECT 77.543 91.669 78.923 91.72 ;
      RECT 77.589 91.623 78.969 91.674 ;
      RECT 77.635 91.577 79.015 91.628 ;
      RECT 77.681 91.531 79.061 91.582 ;
      RECT 77.727 91.485 79.107 91.536 ;
      RECT 77.773 91.439 79.153 91.49 ;
      RECT 77.819 91.393 79.199 91.444 ;
      RECT 77.865 91.347 79.245 91.398 ;
      RECT 77.911 91.301 79.291 91.352 ;
      RECT 77.957 91.255 79.337 91.306 ;
      RECT 78.003 91.209 79.383 91.26 ;
      RECT 78.049 91.163 79.429 91.214 ;
      RECT 78.095 91.117 79.475 91.168 ;
      RECT 78.141 91.071 79.521 91.122 ;
      RECT 78.187 91.025 79.567 91.076 ;
      RECT 78.233 90.979 79.613 91.03 ;
      RECT 78.279 90.933 79.659 90.984 ;
      RECT 78.325 90.887 79.705 90.938 ;
      RECT 78.371 90.841 79.751 90.892 ;
      RECT 78.417 90.795 79.797 90.846 ;
      RECT 78.463 90.749 79.843 90.8 ;
      RECT 78.509 90.703 79.889 90.754 ;
      RECT 78.555 90.657 79.935 90.708 ;
      RECT 78.601 90.611 79.981 90.662 ;
      RECT 78.647 90.565 80.027 90.616 ;
      RECT 78.693 90.519 80.073 90.57 ;
      RECT 78.739 90.473 80.119 90.524 ;
      RECT 78.785 90.427 80.165 90.478 ;
      RECT 78.831 90.381 80.211 90.432 ;
      RECT 78.877 90.335 80.257 90.386 ;
      RECT 78.923 90.289 80.303 90.34 ;
      RECT 78.969 90.243 80.349 90.294 ;
      RECT 79.015 90.197 80.395 90.248 ;
      RECT 79.061 90.151 80.441 90.202 ;
      RECT 79.107 90.105 80.487 90.156 ;
      RECT 79.153 90.059 80.533 90.11 ;
      RECT 79.199 90.013 80.579 90.064 ;
      RECT 79.245 89.967 80.625 90.018 ;
      RECT 79.291 89.921 80.671 89.972 ;
      RECT 79.337 89.875 80.717 89.926 ;
      RECT 79.383 89.829 80.763 89.88 ;
      RECT 79.429 89.783 80.809 89.834 ;
      RECT 79.475 89.737 80.855 89.788 ;
      RECT 79.521 89.691 80.901 89.742 ;
      RECT 79.567 89.645 80.947 89.696 ;
      RECT 79.613 89.599 80.993 89.65 ;
      RECT 79.659 89.553 81.039 89.604 ;
      RECT 79.705 89.507 81.085 89.558 ;
      RECT 79.751 89.461 81.131 89.512 ;
      RECT 79.797 89.415 81.177 89.466 ;
      RECT 79.843 89.369 81.223 89.42 ;
      RECT 79.889 89.323 81.269 89.374 ;
      RECT 79.935 89.277 81.315 89.328 ;
      RECT 79.981 89.231 81.361 89.282 ;
      RECT 80.027 89.185 81.407 89.236 ;
      RECT 80.073 89.139 81.453 89.19 ;
      RECT 80.119 89.093 81.499 89.144 ;
      RECT 80.165 89.047 81.545 89.098 ;
      RECT 80.211 89.001 81.591 89.052 ;
      RECT 80.257 88.955 81.637 89.006 ;
      RECT 80.303 88.909 81.683 88.96 ;
      RECT 80.349 88.863 81.729 88.914 ;
      RECT 80.395 88.817 81.775 88.868 ;
      RECT 80.441 88.771 81.821 88.822 ;
      RECT 80.487 88.725 81.867 88.776 ;
      RECT 80.533 88.679 81.913 88.73 ;
      RECT 80.579 88.633 81.959 88.684 ;
      RECT 80.625 88.587 82.005 88.638 ;
      RECT 80.671 88.541 82.051 88.592 ;
      RECT 80.717 88.495 82.097 88.546 ;
      RECT 80.763 88.449 82.143 88.5 ;
      RECT 80.809 88.403 82.189 88.454 ;
      RECT 80.855 88.357 82.235 88.408 ;
      RECT 80.901 88.311 82.281 88.362 ;
      RECT 80.947 88.265 82.327 88.316 ;
      RECT 80.993 88.219 82.373 88.27 ;
      RECT 81.039 88.173 82.419 88.224 ;
      RECT 81.085 88.127 82.465 88.178 ;
      RECT 81.131 88.081 82.511 88.132 ;
      RECT 81.177 88.035 82.557 88.086 ;
      RECT 81.223 87.989 82.603 88.04 ;
      RECT 81.269 87.943 82.649 87.994 ;
      RECT 81.315 87.897 82.695 87.948 ;
      RECT 81.361 87.851 82.741 87.902 ;
      RECT 81.407 87.805 82.787 87.856 ;
      RECT 81.453 87.759 82.833 87.81 ;
      RECT 81.499 87.713 82.879 87.764 ;
      RECT 81.545 87.667 82.925 87.718 ;
      RECT 81.591 87.621 82.971 87.672 ;
      RECT 81.637 87.575 83.017 87.626 ;
      RECT 81.683 87.529 83.063 87.58 ;
      RECT 81.729 87.483 83.109 87.534 ;
      RECT 81.775 87.437 83.155 87.488 ;
      RECT 81.821 87.391 83.201 87.442 ;
      RECT 81.867 87.345 83.247 87.396 ;
      RECT 81.913 87.299 83.293 87.35 ;
      RECT 81.959 87.253 83.339 87.304 ;
      RECT 82.005 87.207 83.385 87.258 ;
      RECT 82.051 87.161 83.431 87.212 ;
      RECT 82.097 87.115 83.477 87.166 ;
      RECT 82.143 87.069 83.523 87.12 ;
      RECT 82.189 87.023 83.569 87.074 ;
      RECT 82.235 86.977 83.615 87.028 ;
      RECT 82.281 86.931 83.661 86.982 ;
      RECT 82.327 86.885 83.707 86.936 ;
      RECT 82.373 86.839 83.753 86.89 ;
      RECT 82.419 86.793 83.799 86.844 ;
      RECT 82.465 86.747 83.845 86.798 ;
      RECT 82.511 86.701 83.891 86.752 ;
      RECT 82.557 86.655 83.937 86.706 ;
      RECT 82.603 86.609 83.983 86.66 ;
      RECT 82.649 86.563 84.029 86.614 ;
      RECT 82.695 86.517 84.075 86.568 ;
      RECT 82.741 86.471 84.121 86.522 ;
      RECT 82.787 86.425 84.167 86.476 ;
      RECT 82.833 86.379 84.213 86.43 ;
      RECT 82.879 86.333 84.259 86.384 ;
      RECT 82.925 86.287 84.305 86.338 ;
      RECT 82.971 86.241 84.351 86.292 ;
      RECT 83.017 86.195 84.397 86.246 ;
      RECT 83.063 86.149 84.443 86.2 ;
      RECT 83.109 86.103 84.489 86.154 ;
      RECT 83.155 86.057 84.535 86.108 ;
      RECT 83.201 86.011 84.581 86.062 ;
      RECT 83.247 85.965 84.627 86.016 ;
      RECT 83.293 85.919 84.673 85.97 ;
      RECT 83.339 85.873 84.719 85.924 ;
      RECT 83.385 85.827 84.765 85.878 ;
      RECT 83.431 85.781 84.811 85.832 ;
      RECT 83.477 85.735 84.857 85.786 ;
      RECT 83.523 85.689 84.903 85.74 ;
      RECT 83.569 85.643 84.949 85.694 ;
      RECT 83.615 85.597 84.995 85.648 ;
      RECT 83.661 85.551 85.041 85.602 ;
      RECT 83.707 85.505 85.087 85.556 ;
      RECT 83.753 85.459 85.133 85.51 ;
      RECT 83.799 85.413 85.179 85.464 ;
      RECT 83.845 85.367 85.225 85.418 ;
      RECT 83.891 85.321 85.271 85.372 ;
      RECT 83.937 85.275 85.317 85.326 ;
      RECT 83.983 85.229 85.363 85.28 ;
      RECT 84.029 85.183 85.409 85.234 ;
      RECT 84.075 85.137 85.455 85.188 ;
      RECT 84.121 85.091 85.501 85.142 ;
      RECT 84.167 85.045 85.547 85.096 ;
      RECT 84.213 84.999 85.593 85.05 ;
      RECT 84.259 84.953 85.639 85.004 ;
      RECT 84.305 84.907 85.685 84.958 ;
      RECT 84.351 84.861 85.731 84.912 ;
      RECT 84.397 84.815 85.777 84.866 ;
      RECT 84.443 84.769 85.823 84.82 ;
      RECT 84.489 84.723 85.869 84.774 ;
      RECT 84.535 84.677 85.915 84.728 ;
      RECT 84.581 84.631 85.961 84.682 ;
      RECT 84.627 84.585 86.007 84.636 ;
      RECT 84.673 84.539 86.053 84.59 ;
      RECT 84.719 84.493 86.099 84.544 ;
      RECT 84.765 84.447 86.145 84.498 ;
      RECT 84.811 84.401 86.191 84.452 ;
      RECT 84.857 84.355 86.237 84.406 ;
      RECT 84.903 84.309 86.283 84.36 ;
      RECT 84.949 84.263 86.329 84.314 ;
      RECT 84.995 84.217 86.375 84.268 ;
      RECT 85.041 84.171 86.421 84.222 ;
      RECT 85.087 84.125 86.467 84.176 ;
      RECT 85.133 84.079 86.513 84.13 ;
      RECT 85.179 84.033 86.559 84.084 ;
      RECT 85.225 83.987 86.605 84.038 ;
      RECT 85.271 83.941 86.651 83.992 ;
      RECT 85.317 83.895 86.697 83.946 ;
      RECT 85.363 83.849 86.743 83.9 ;
      RECT 85.409 83.803 86.789 83.854 ;
      RECT 85.455 83.757 86.835 83.808 ;
      RECT 85.501 83.711 86.881 83.762 ;
      RECT 85.547 83.665 86.927 83.716 ;
      RECT 85.593 83.619 86.973 83.67 ;
      RECT 85.639 83.573 87.019 83.624 ;
      RECT 85.685 83.527 87.065 83.578 ;
      RECT 85.731 83.481 87.111 83.532 ;
      RECT 85.777 83.435 87.157 83.486 ;
      RECT 85.823 83.389 87.203 83.44 ;
      RECT 85.869 83.343 87.249 83.394 ;
      RECT 85.915 83.297 87.295 83.348 ;
      RECT 85.961 83.251 87.341 83.302 ;
      RECT 86.007 83.205 87.387 83.256 ;
      RECT 86.053 83.159 87.433 83.21 ;
      RECT 86.099 83.113 87.479 83.164 ;
      RECT 86.145 83.067 87.525 83.118 ;
      RECT 86.191 83.021 87.571 83.072 ;
      RECT 86.237 82.975 87.617 83.026 ;
      RECT 86.283 82.929 87.663 82.98 ;
      RECT 86.329 82.883 87.709 82.934 ;
      RECT 86.375 82.837 87.755 82.888 ;
      RECT 86.421 82.791 87.801 82.842 ;
      RECT 86.467 82.745 87.847 82.796 ;
      RECT 86.513 82.699 87.893 82.75 ;
      RECT 86.559 82.653 87.939 82.704 ;
      RECT 86.605 82.607 87.985 82.658 ;
      RECT 86.651 82.561 88.031 82.612 ;
      RECT 86.697 82.515 88.077 82.566 ;
      RECT 86.743 82.469 88.123 82.52 ;
      RECT 86.789 82.423 88.169 82.474 ;
      RECT 86.835 82.377 88.215 82.428 ;
      RECT 86.881 82.331 88.261 82.382 ;
      RECT 86.927 82.285 88.307 82.336 ;
      RECT 86.973 82.239 88.353 82.29 ;
      RECT 87.019 82.193 88.399 82.244 ;
      RECT 87.065 82.147 88.445 82.198 ;
      RECT 87.111 82.101 88.491 82.152 ;
      RECT 87.157 82.055 88.537 82.106 ;
      RECT 87.203 82.009 88.583 82.06 ;
      RECT 88.537 80.697 88.583 82.06 ;
      RECT 87.249 81.963 88.629 82.014 ;
      RECT 87.295 81.917 88.675 81.968 ;
      RECT 87.341 81.871 88.721 81.922 ;
      RECT 87.387 81.825 88.767 81.876 ;
      RECT 87.433 81.779 88.813 81.83 ;
      RECT 87.479 81.733 88.859 81.784 ;
      RECT 87.525 81.687 88.905 81.738 ;
      RECT 87.571 81.641 88.951 81.692 ;
      RECT 87.617 81.595 88.997 81.646 ;
      RECT 87.663 81.549 89.043 81.6 ;
      RECT 87.709 81.503 89.089 81.554 ;
      RECT 87.755 81.457 89.135 81.508 ;
      RECT 87.801 81.411 89.181 81.462 ;
      RECT 87.847 81.365 89.227 81.416 ;
      RECT 87.893 81.319 89.273 81.37 ;
      RECT 87.939 81.273 89.319 81.324 ;
      RECT 87.939 81.273 89.325 81.298 ;
      RECT 87.985 81.227 89.371 81.272 ;
      RECT 88.031 81.181 89.417 81.226 ;
      RECT 88.077 81.135 89.463 81.18 ;
      RECT 88.123 81.089 89.509 81.134 ;
      RECT 88.169 81.043 89.555 81.088 ;
      RECT 88.215 80.997 89.601 81.042 ;
      RECT 88.261 80.951 89.647 80.996 ;
      RECT 88.307 80.905 89.693 80.95 ;
      RECT 88.353 80.859 89.739 80.904 ;
      RECT 88.399 80.813 89.785 80.858 ;
      RECT 88.445 80.767 89.831 80.812 ;
      RECT 88.491 80.721 89.877 80.766 ;
      RECT 88.54 80.672 89.923 80.72 ;
      RECT 89.874 79.338 89.923 80.72 ;
      RECT 88.586 80.626 89.969 80.674 ;
      RECT 89.92 79.292 89.969 80.674 ;
      RECT 88.632 80.58 90.015 80.628 ;
      RECT 89.966 79.246 90.015 80.628 ;
      RECT 88.678 80.534 90.061 80.582 ;
      RECT 90.012 79.2 90.061 80.582 ;
      RECT 88.724 80.488 90.107 80.536 ;
      RECT 90.058 79.154 90.107 80.536 ;
      RECT 88.77 80.442 90.153 80.49 ;
      RECT 90.104 79.108 90.153 80.49 ;
      RECT 88.816 80.396 90.199 80.444 ;
      RECT 90.15 79.062 90.199 80.444 ;
      RECT 88.862 80.35 90.245 80.398 ;
      RECT 90.196 79.016 90.245 80.398 ;
      RECT 88.908 80.304 90.291 80.352 ;
      RECT 90.242 78.97 90.291 80.352 ;
      RECT 88.954 80.258 90.337 80.306 ;
      RECT 90.288 78.924 90.337 80.306 ;
      RECT 89 80.212 90.383 80.26 ;
      RECT 90.334 78.878 90.383 80.26 ;
      RECT 89.046 80.166 90.429 80.214 ;
      RECT 90.38 78.832 90.429 80.214 ;
      RECT 89.092 80.12 90.475 80.168 ;
      RECT 90.426 78.786 90.475 80.168 ;
      RECT 89.138 80.074 90.521 80.122 ;
      RECT 90.472 78.74 90.521 80.122 ;
      RECT 89.184 80.028 90.567 80.076 ;
      RECT 90.518 78.694 90.567 80.076 ;
      RECT 89.23 79.982 90.613 80.03 ;
      RECT 90.564 78.648 90.613 80.03 ;
      RECT 89.276 79.936 90.659 79.984 ;
      RECT 90.61 78.602 90.659 79.984 ;
      RECT 89.322 79.89 90.705 79.938 ;
      RECT 90.656 78.556 90.705 79.938 ;
      RECT 89.368 79.844 90.751 79.892 ;
      RECT 90.702 78.51 90.751 79.892 ;
      RECT 89.414 79.798 90.797 79.846 ;
      RECT 90.748 78.464 90.797 79.846 ;
      RECT 89.46 79.752 90.843 79.8 ;
      RECT 90.794 78.418 90.843 79.8 ;
      RECT 89.506 79.706 90.889 79.754 ;
      RECT 90.84 78.372 90.889 79.754 ;
      RECT 89.552 79.66 90.935 79.708 ;
      RECT 90.886 78.326 90.935 79.708 ;
      RECT 89.598 79.614 90.981 79.662 ;
      RECT 90.932 78.28 90.981 79.662 ;
      RECT 89.644 79.568 91.027 79.616 ;
      RECT 90.978 78.234 91.027 79.616 ;
      RECT 89.69 79.522 91.073 79.57 ;
      RECT 91.024 78.188 91.073 79.57 ;
      RECT 89.736 79.476 91.119 79.524 ;
      RECT 91.07 78.142 91.119 79.524 ;
      RECT 89.782 79.43 91.165 79.478 ;
      RECT 91.116 78.096 91.165 79.478 ;
      RECT 89.828 79.384 91.211 79.432 ;
      RECT 91.162 78.05 91.211 79.432 ;
      RECT 91.208 78.004 91.257 79.386 ;
      RECT 91.254 77.958 91.303 79.34 ;
      RECT 91.3 77.912 91.349 79.294 ;
      RECT 91.346 77.866 91.395 79.248 ;
      RECT 91.392 77.82 91.441 79.202 ;
      RECT 91.438 77.774 91.487 79.156 ;
      RECT 91.484 77.728 91.533 79.11 ;
      RECT 91.53 77.682 91.579 79.064 ;
      RECT 91.576 77.636 91.625 79.018 ;
      RECT 91.622 77.59 91.671 78.972 ;
      RECT 91.668 77.544 91.717 78.926 ;
      RECT 91.714 77.498 91.763 78.88 ;
      RECT 91.76 77.452 91.809 78.834 ;
      RECT 91.806 77.406 91.855 78.788 ;
      RECT 91.852 77.36 91.901 78.742 ;
      RECT 91.898 77.314 91.947 78.696 ;
      RECT 91.944 77.268 91.993 78.65 ;
      RECT 91.99 77.222 92.039 78.604 ;
      RECT 92.036 77.187 92.085 78.558 ;
      RECT 92.06 77.175 92.131 78.512 ;
      RECT 92.06 77.175 92.177 78.466 ;
      RECT 92.06 77.175 92.223 78.42 ;
      RECT 92.06 77.175 92.269 78.374 ;
      RECT 90.886 78.326 92.295 78.338 ;
      RECT 92.06 77.175 110 78.325 ;
      RECT 89.675 97.182 90.825 110 ;
      RECT 89.675 97.182 90.871 99.352 ;
      RECT 89.675 97.182 90.917 99.306 ;
      RECT 89.675 97.182 90.963 99.26 ;
      RECT 89.675 97.182 91.009 99.214 ;
      RECT 89.675 97.182 91.055 99.168 ;
      RECT 89.675 97.182 91.101 99.122 ;
      RECT 89.675 97.182 91.147 99.076 ;
      RECT 89.675 97.182 91.193 99.03 ;
      RECT 89.675 97.182 91.239 98.984 ;
      RECT 89.675 97.182 91.285 98.938 ;
      RECT 89.675 97.182 91.331 98.892 ;
      RECT 89.675 97.182 91.377 98.846 ;
      RECT 89.675 97.182 91.423 98.8 ;
      RECT 89.675 97.182 91.469 98.754 ;
      RECT 89.675 97.182 91.515 98.708 ;
      RECT 89.675 97.182 91.561 98.662 ;
      RECT 89.675 97.182 91.607 98.616 ;
      RECT 89.675 97.182 91.653 98.57 ;
      RECT 89.675 97.182 91.699 98.524 ;
      RECT 89.675 97.182 91.745 98.478 ;
      RECT 89.675 97.182 91.791 98.432 ;
      RECT 89.675 97.182 91.837 98.386 ;
      RECT 89.675 97.182 91.883 98.34 ;
      RECT 89.675 97.182 91.929 98.294 ;
      RECT 89.675 97.182 91.975 98.248 ;
      RECT 89.675 97.182 92.021 98.202 ;
      RECT 89.675 97.182 92.067 98.156 ;
      RECT 89.675 97.182 92.113 98.11 ;
      RECT 89.675 97.182 92.159 98.064 ;
      RECT 89.675 97.182 92.205 98.018 ;
      RECT 89.675 97.182 92.251 97.972 ;
      RECT 89.675 97.182 92.297 97.926 ;
      RECT 89.675 97.182 92.343 97.88 ;
      RECT 89.675 97.182 92.389 97.834 ;
      RECT 89.675 97.182 92.435 97.788 ;
      RECT 89.675 97.182 92.481 97.742 ;
      RECT 89.675 97.182 92.527 97.696 ;
      RECT 89.675 97.182 92.573 97.65 ;
      RECT 89.675 97.182 92.619 97.604 ;
      RECT 89.675 97.182 92.665 97.558 ;
      RECT 89.675 97.182 92.711 97.512 ;
      RECT 89.675 97.182 92.757 97.466 ;
      RECT 89.675 97.182 92.803 97.42 ;
      RECT 89.675 97.182 92.849 97.374 ;
      RECT 89.675 97.182 92.895 97.328 ;
      RECT 89.675 97.182 92.941 97.282 ;
      RECT 89.721 97.136 93.033 97.19 ;
      RECT 92.967 93.89 93.033 97.19 ;
      RECT 89.767 97.09 93.079 97.144 ;
      RECT 93.013 93.844 93.079 97.144 ;
      RECT 89.813 97.044 93.125 97.098 ;
      RECT 93.059 93.798 93.125 97.098 ;
      RECT 89.859 96.998 93.171 97.052 ;
      RECT 93.105 93.752 93.171 97.052 ;
      RECT 89.905 96.952 93.217 97.006 ;
      RECT 93.151 93.706 93.217 97.006 ;
      RECT 89.951 96.906 93.263 96.96 ;
      RECT 93.197 93.66 93.263 96.96 ;
      RECT 89.997 96.86 93.309 96.914 ;
      RECT 93.243 93.614 93.309 96.914 ;
      RECT 90.043 96.814 93.355 96.868 ;
      RECT 93.289 93.568 93.355 96.868 ;
      RECT 90.089 96.768 93.401 96.822 ;
      RECT 93.335 93.522 93.401 96.822 ;
      RECT 90.135 96.722 93.447 96.776 ;
      RECT 93.381 93.476 93.447 96.776 ;
      RECT 90.181 96.676 93.493 96.73 ;
      RECT 93.427 93.43 93.493 96.73 ;
      RECT 90.227 96.63 93.539 96.684 ;
      RECT 93.473 93.384 93.539 96.684 ;
      RECT 90.273 96.584 93.585 96.638 ;
      RECT 93.519 93.338 93.585 96.638 ;
      RECT 90.319 96.538 93.631 96.592 ;
      RECT 93.565 93.292 93.631 96.592 ;
      RECT 90.365 96.492 93.677 96.546 ;
      RECT 93.611 93.246 93.677 96.546 ;
      RECT 90.411 96.446 93.723 96.5 ;
      RECT 93.657 93.2 93.723 96.5 ;
      RECT 90.457 96.4 93.769 96.454 ;
      RECT 93.703 93.154 93.769 96.454 ;
      RECT 90.503 96.354 93.815 96.408 ;
      RECT 93.749 93.108 93.815 96.408 ;
      RECT 90.549 96.308 93.861 96.362 ;
      RECT 93.795 93.062 93.861 96.362 ;
      RECT 90.595 96.262 93.907 96.316 ;
      RECT 93.841 93.016 93.907 96.316 ;
      RECT 90.641 96.216 93.953 96.27 ;
      RECT 93.887 92.97 93.953 96.27 ;
      RECT 90.687 96.17 93.999 96.224 ;
      RECT 93.933 92.924 93.999 96.224 ;
      RECT 90.733 96.124 94.045 96.178 ;
      RECT 93.979 92.878 94.045 96.178 ;
      RECT 90.779 96.078 94.091 96.132 ;
      RECT 94.025 92.832 94.091 96.132 ;
      RECT 90.825 96.032 94.137 96.086 ;
      RECT 94.071 92.786 94.137 96.086 ;
      RECT 90.871 95.986 94.183 96.04 ;
      RECT 94.117 92.74 94.183 96.04 ;
      RECT 90.917 95.94 94.229 95.994 ;
      RECT 94.163 92.694 94.229 95.994 ;
      RECT 90.963 95.894 94.275 95.948 ;
      RECT 94.209 92.648 94.275 95.948 ;
      RECT 91.009 95.848 94.321 95.902 ;
      RECT 94.255 92.602 94.321 95.902 ;
      RECT 91.055 95.802 94.367 95.856 ;
      RECT 94.301 92.556 94.367 95.856 ;
      RECT 91.101 95.756 94.413 95.81 ;
      RECT 94.347 92.51 94.413 95.81 ;
      RECT 91.147 95.71 94.459 95.764 ;
      RECT 94.393 92.464 94.459 95.764 ;
      RECT 91.193 95.664 94.505 95.718 ;
      RECT 94.439 92.418 94.505 95.718 ;
      RECT 91.239 95.618 94.551 95.672 ;
      RECT 94.485 92.372 94.551 95.672 ;
      RECT 91.285 95.572 94.597 95.626 ;
      RECT 94.531 92.326 94.597 95.626 ;
      RECT 91.331 95.526 94.643 95.58 ;
      RECT 94.577 92.28 94.643 95.58 ;
      RECT 91.377 95.48 94.689 95.534 ;
      RECT 94.623 92.234 94.689 95.534 ;
      RECT 91.423 95.434 94.735 95.488 ;
      RECT 94.669 92.188 94.735 95.488 ;
      RECT 91.469 95.388 94.781 95.442 ;
      RECT 94.715 92.142 94.781 95.442 ;
      RECT 91.515 95.342 94.827 95.396 ;
      RECT 94.761 92.096 94.827 95.396 ;
      RECT 91.561 95.296 94.873 95.35 ;
      RECT 94.807 92.05 94.873 95.35 ;
      RECT 91.607 95.25 94.919 95.304 ;
      RECT 94.853 92.004 94.919 95.304 ;
      RECT 91.653 95.204 94.965 95.258 ;
      RECT 94.899 91.958 94.965 95.258 ;
      RECT 91.699 95.158 95.011 95.212 ;
      RECT 94.945 91.912 95.011 95.212 ;
      RECT 91.745 95.112 95.057 95.166 ;
      RECT 94.991 91.866 95.057 95.166 ;
      RECT 91.791 95.066 95.103 95.12 ;
      RECT 95.037 91.82 95.103 95.12 ;
      RECT 91.837 95.02 95.149 95.074 ;
      RECT 95.083 91.774 95.149 95.074 ;
      RECT 91.883 94.974 95.195 95.028 ;
      RECT 95.129 91.728 95.195 95.028 ;
      RECT 91.929 94.928 95.241 94.982 ;
      RECT 95.175 91.682 95.241 94.982 ;
      RECT 91.975 94.882 95.287 94.936 ;
      RECT 95.221 91.636 95.287 94.936 ;
      RECT 92.021 94.836 95.333 94.89 ;
      RECT 95.267 91.59 95.333 94.89 ;
      RECT 92.067 94.79 95.379 94.844 ;
      RECT 95.313 91.544 95.379 94.844 ;
      RECT 92.113 94.744 95.425 94.798 ;
      RECT 95.359 91.498 95.425 94.798 ;
      RECT 92.159 94.698 95.471 94.752 ;
      RECT 95.405 91.452 95.471 94.752 ;
      RECT 92.205 94.652 95.517 94.706 ;
      RECT 95.451 91.406 95.517 94.706 ;
      RECT 92.251 94.606 95.563 94.66 ;
      RECT 95.497 91.36 95.563 94.66 ;
      RECT 92.297 94.56 95.609 94.614 ;
      RECT 95.543 91.314 95.609 94.614 ;
      RECT 92.343 94.514 95.655 94.568 ;
      RECT 95.589 91.268 95.655 94.568 ;
      RECT 92.389 94.468 95.701 94.522 ;
      RECT 95.635 91.222 95.701 94.522 ;
      RECT 92.435 94.422 95.747 94.476 ;
      RECT 95.681 91.176 95.747 94.476 ;
      RECT 92.481 94.376 95.793 94.43 ;
      RECT 95.727 91.13 95.793 94.43 ;
      RECT 92.527 94.33 95.839 94.384 ;
      RECT 95.773 91.084 95.839 94.384 ;
      RECT 92.573 94.284 95.885 94.338 ;
      RECT 95.819 91.038 95.885 94.338 ;
      RECT 92.619 94.248 95.931 94.292 ;
      RECT 95.865 90.992 95.931 94.292 ;
      RECT 92.645 94.212 95.931 94.292 ;
      RECT 92.921 93.936 92.987 97.236 ;
      RECT 92.691 94.166 95.977 94.246 ;
      RECT 95.911 90.946 95.977 94.246 ;
      RECT 92.737 94.12 96.023 94.2 ;
      RECT 95.957 90.9 96.023 94.2 ;
      RECT 92.783 94.074 96.069 94.154 ;
      RECT 96.003 90.854 96.069 94.154 ;
      RECT 92.829 94.028 96.115 94.108 ;
      RECT 96.049 90.808 96.115 94.108 ;
      RECT 92.875 93.982 96.161 94.062 ;
      RECT 96.095 90.762 96.161 94.062 ;
      RECT 96.141 90.716 96.207 94.016 ;
      RECT 96.187 90.67 96.253 93.97 ;
      RECT 96.233 90.624 96.299 93.924 ;
      RECT 96.279 90.578 96.345 93.878 ;
      RECT 96.325 90.532 96.391 93.832 ;
      RECT 96.371 90.486 96.437 93.786 ;
      RECT 96.417 90.44 96.483 93.74 ;
      RECT 96.463 90.394 96.529 93.694 ;
      RECT 96.509 90.348 96.575 93.648 ;
      RECT 96.555 90.302 96.621 93.602 ;
      RECT 96.601 90.256 96.667 93.556 ;
      RECT 96.647 90.21 96.713 93.51 ;
      RECT 96.693 90.164 96.759 93.464 ;
      RECT 96.739 90.118 96.805 93.418 ;
      RECT 96.785 90.072 96.851 93.372 ;
      RECT 96.831 90.026 96.897 93.326 ;
      RECT 96.877 89.98 96.943 93.28 ;
      RECT 96.923 89.934 96.989 93.234 ;
      RECT 96.969 89.888 97.035 93.188 ;
      RECT 97.015 89.842 97.081 93.142 ;
      RECT 97.061 89.796 97.127 93.096 ;
      RECT 97.107 89.75 97.173 93.05 ;
      RECT 97.199 89.678 97.219 93.004 ;
      RECT 97.205 89.675 97.265 92.958 ;
      RECT 97.153 89.704 97.219 93.004 ;
      RECT 97.205 89.675 97.311 92.912 ;
      RECT 97.205 89.675 97.357 92.866 ;
      RECT 97.205 89.675 97.403 92.82 ;
      RECT 97.205 89.675 97.449 92.774 ;
      RECT 97.205 89.675 97.495 92.728 ;
      RECT 97.205 89.675 97.541 92.682 ;
      RECT 97.205 89.675 97.587 92.636 ;
      RECT 97.205 89.675 97.633 92.59 ;
      RECT 97.205 89.675 97.679 92.544 ;
      RECT 97.205 89.675 97.725 92.498 ;
      RECT 97.205 89.675 97.771 92.452 ;
      RECT 94.485 92.372 97.817 92.406 ;
      RECT 97.205 89.675 97.825 92.379 ;
      RECT 97.205 89.675 97.871 92.352 ;
      RECT 97.205 89.675 97.917 92.306 ;
      RECT 97.205 89.675 97.963 92.26 ;
      RECT 97.205 89.675 98.009 92.214 ;
      RECT 97.205 89.675 98.055 92.168 ;
      RECT 97.205 89.675 98.101 92.122 ;
      RECT 97.205 89.675 98.147 92.076 ;
      RECT 97.205 89.675 98.193 92.03 ;
      RECT 97.205 89.675 98.239 91.984 ;
      RECT 97.205 89.675 98.285 91.938 ;
      RECT 97.205 89.675 98.331 91.892 ;
      RECT 97.205 89.675 98.377 91.846 ;
      RECT 97.205 89.675 98.423 91.8 ;
      RECT 97.205 89.675 98.469 91.754 ;
      RECT 97.205 89.675 98.515 91.708 ;
      RECT 97.205 89.675 98.561 91.662 ;
      RECT 97.205 89.675 98.607 91.616 ;
      RECT 97.205 89.675 98.653 91.57 ;
      RECT 97.205 89.675 98.699 91.524 ;
      RECT 97.205 89.675 98.745 91.478 ;
      RECT 97.205 89.675 98.791 91.432 ;
      RECT 97.205 89.675 98.837 91.386 ;
      RECT 97.205 89.675 98.883 91.34 ;
      RECT 97.205 89.675 98.929 91.294 ;
      RECT 97.205 89.675 98.975 91.248 ;
      RECT 97.205 89.675 99.021 91.202 ;
      RECT 97.205 89.675 99.067 91.156 ;
      RECT 97.205 89.675 99.113 91.11 ;
      RECT 97.205 89.675 99.159 91.064 ;
      RECT 97.205 89.675 99.205 91.018 ;
      RECT 97.205 89.675 99.251 90.972 ;
      RECT 97.205 89.675 99.297 90.926 ;
      RECT 97.205 89.675 99.343 90.88 ;
      RECT 96.049 90.808 99.375 90.841 ;
      RECT 97.205 89.675 110 90.825 ;
      RECT 98.175 102.602 99.325 110 ;
      RECT 98.175 102.602 99.371 103.642 ;
      RECT 98.175 102.602 99.417 103.596 ;
      RECT 98.175 102.602 99.463 103.55 ;
      RECT 98.175 102.602 99.509 103.504 ;
      RECT 98.175 102.602 99.555 103.458 ;
      RECT 98.175 102.602 99.601 103.412 ;
      RECT 98.175 102.602 99.647 103.366 ;
      RECT 98.175 102.602 99.693 103.32 ;
      RECT 98.175 102.602 99.739 103.274 ;
      RECT 98.175 102.602 99.785 103.228 ;
      RECT 98.175 102.602 99.831 103.182 ;
      RECT 98.175 102.602 99.877 103.136 ;
      RECT 98.175 102.602 99.923 103.09 ;
      RECT 98.175 102.602 99.969 103.044 ;
      RECT 98.175 102.602 100.015 102.998 ;
      RECT 98.175 102.602 100.061 102.952 ;
      RECT 98.175 102.602 100.107 102.906 ;
      RECT 98.175 102.602 100.153 102.86 ;
      RECT 98.175 102.602 100.199 102.814 ;
      RECT 98.175 102.602 100.245 102.768 ;
      RECT 98.175 102.602 100.291 102.722 ;
      RECT 98.175 102.602 100.337 102.676 ;
      RECT 98.221 102.556 100.383 102.63 ;
      RECT 100.323 100.454 100.383 102.63 ;
      RECT 98.267 102.51 100.429 102.584 ;
      RECT 100.369 100.408 100.429 102.584 ;
      RECT 98.313 102.464 100.475 102.538 ;
      RECT 100.415 100.362 100.475 102.538 ;
      RECT 98.359 102.418 100.521 102.492 ;
      RECT 100.461 100.316 100.521 102.492 ;
      RECT 98.405 102.372 100.567 102.446 ;
      RECT 100.507 100.27 100.567 102.446 ;
      RECT 98.451 102.326 100.613 102.4 ;
      RECT 100.553 100.224 100.613 102.4 ;
      RECT 98.497 102.28 100.659 102.354 ;
      RECT 100.599 100.178 100.659 102.354 ;
      RECT 98.543 102.234 100.705 102.308 ;
      RECT 100.645 100.132 100.705 102.308 ;
      RECT 98.589 102.188 100.751 102.262 ;
      RECT 100.691 100.086 100.751 102.262 ;
      RECT 98.635 102.142 100.797 102.216 ;
      RECT 100.737 100.04 100.797 102.216 ;
      RECT 98.681 102.096 100.843 102.17 ;
      RECT 100.783 99.994 100.843 102.17 ;
      RECT 98.727 102.05 100.889 102.124 ;
      RECT 100.829 99.948 100.889 102.124 ;
      RECT 98.773 102.004 100.935 102.078 ;
      RECT 100.875 99.902 100.935 102.078 ;
      RECT 98.819 101.958 100.981 102.032 ;
      RECT 100.921 99.856 100.981 102.032 ;
      RECT 98.865 101.912 101.027 101.986 ;
      RECT 100.967 99.81 101.027 101.986 ;
      RECT 98.911 101.866 101.073 101.94 ;
      RECT 101.013 99.764 101.073 101.94 ;
      RECT 98.957 101.82 101.119 101.894 ;
      RECT 101.059 99.718 101.119 101.894 ;
      RECT 99.003 101.774 101.165 101.848 ;
      RECT 101.105 99.672 101.165 101.848 ;
      RECT 99.049 101.728 101.211 101.802 ;
      RECT 101.151 99.626 101.211 101.802 ;
      RECT 99.095 101.682 101.257 101.756 ;
      RECT 101.197 99.58 101.257 101.756 ;
      RECT 99.141 101.636 101.303 101.71 ;
      RECT 101.243 99.534 101.303 101.71 ;
      RECT 99.187 101.59 101.349 101.664 ;
      RECT 101.289 99.488 101.349 101.664 ;
      RECT 99.233 101.544 101.395 101.618 ;
      RECT 101.335 99.442 101.395 101.618 ;
      RECT 99.279 101.498 101.441 101.572 ;
      RECT 101.381 99.396 101.441 101.572 ;
      RECT 99.325 101.452 101.487 101.526 ;
      RECT 101.427 99.35 101.487 101.526 ;
      RECT 99.371 101.406 101.533 101.48 ;
      RECT 101.473 99.304 101.533 101.48 ;
      RECT 99.417 101.36 101.579 101.434 ;
      RECT 101.519 99.258 101.579 101.434 ;
      RECT 99.463 101.314 101.625 101.388 ;
      RECT 101.565 99.212 101.625 101.388 ;
      RECT 99.509 101.268 101.671 101.342 ;
      RECT 101.611 99.166 101.671 101.342 ;
      RECT 99.555 101.222 101.717 101.296 ;
      RECT 101.657 99.12 101.717 101.296 ;
      RECT 99.601 101.176 101.763 101.25 ;
      RECT 101.703 99.074 101.763 101.25 ;
      RECT 99.647 101.13 101.809 101.204 ;
      RECT 101.749 99.028 101.809 101.204 ;
      RECT 99.693 101.091 101.855 101.158 ;
      RECT 101.795 98.982 101.855 101.158 ;
      RECT 99.725 101.052 101.901 101.112 ;
      RECT 101.841 98.936 101.901 101.112 ;
      RECT 99.771 101.006 101.947 101.066 ;
      RECT 101.887 98.89 101.947 101.066 ;
      RECT 99.817 100.96 101.993 101.02 ;
      RECT 101.933 98.844 101.993 101.02 ;
      RECT 99.863 100.914 102.039 100.974 ;
      RECT 101.979 98.798 102.039 100.974 ;
      RECT 99.909 100.868 102.085 100.928 ;
      RECT 102.025 98.752 102.085 100.928 ;
      RECT 99.955 100.822 102.131 100.882 ;
      RECT 102.071 98.706 102.131 100.882 ;
      RECT 100.001 100.776 102.177 100.836 ;
      RECT 102.117 98.66 102.177 100.836 ;
      RECT 100.047 100.73 102.223 100.79 ;
      RECT 102.163 98.614 102.223 100.79 ;
      RECT 100.093 100.684 102.269 100.744 ;
      RECT 102.209 98.568 102.269 100.744 ;
      RECT 100.139 100.638 102.315 100.698 ;
      RECT 102.255 98.522 102.315 100.698 ;
      RECT 100.185 100.592 102.361 100.652 ;
      RECT 102.301 98.476 102.361 100.652 ;
      RECT 100.231 100.546 102.407 100.606 ;
      RECT 102.347 98.43 102.407 100.606 ;
      RECT 100.277 100.5 102.453 100.56 ;
      RECT 102.393 98.384 102.453 100.56 ;
      RECT 102.439 98.338 102.499 100.514 ;
      RECT 102.485 98.292 102.545 100.468 ;
      RECT 102.531 98.246 102.591 100.422 ;
      RECT 102.577 98.199 102.637 100.376 ;
      RECT 102.623 98.175 102.683 100.33 ;
      RECT 102.623 98.175 102.729 100.284 ;
      RECT 102.623 98.175 102.775 100.238 ;
      RECT 102.623 98.175 102.821 100.192 ;
      RECT 102.623 98.175 102.867 100.146 ;
      RECT 102.623 98.175 102.913 100.1 ;
      RECT 102.623 98.175 102.959 100.054 ;
      RECT 102.623 98.175 103.005 100.008 ;
      RECT 102.623 98.175 103.051 99.962 ;
      RECT 102.623 98.175 103.097 99.916 ;
      RECT 102.623 98.175 103.143 99.87 ;
      RECT 102.623 98.175 103.189 99.824 ;
      RECT 102.623 98.175 103.235 99.778 ;
      RECT 102.623 98.175 103.281 99.732 ;
      RECT 102.623 98.175 103.327 99.686 ;
      RECT 102.623 98.175 103.373 99.64 ;
      RECT 102.623 98.175 103.419 99.594 ;
      RECT 102.623 98.175 103.465 99.548 ;
      RECT 102.623 98.175 103.511 99.502 ;
      RECT 102.623 98.175 103.557 99.456 ;
      RECT 102.623 98.175 103.603 99.41 ;
      RECT 102.623 98.175 103.649 99.364 ;
      RECT 101.473 99.304 103.665 99.333 ;
      RECT 102.623 98.175 110 99.325 ;
      RECT 107.675 108.902 110 110 ;
      RECT 108.925 107.675 110 110 ;
      RECT 107.721 108.856 110 110 ;
      RECT 108.917 107.679 110 110 ;
      RECT 107.767 108.81 110 110 ;
      RECT 108.871 107.706 110 110 ;
      RECT 107.813 108.764 110 110 ;
      RECT 108.825 107.752 110 110 ;
      RECT 107.859 108.718 110 110 ;
      RECT 108.779 107.798 110 110 ;
      RECT 107.905 108.672 110 110 ;
      RECT 108.733 107.844 110 110 ;
      RECT 107.951 108.626 110 110 ;
      RECT 108.687 107.89 110 110 ;
      RECT 107.997 108.58 110 110 ;
      RECT 108.641 107.936 110 110 ;
      RECT 108.043 108.534 110 110 ;
      RECT 108.595 107.982 110 110 ;
      RECT 108.089 108.488 110 110 ;
      RECT 108.549 108.028 110 110 ;
      RECT 108.135 108.442 110 110 ;
      RECT 108.503 108.074 110 110 ;
      RECT 108.181 108.396 110 110 ;
      RECT 108.457 108.12 110 110 ;
      RECT 108.227 108.35 110 110 ;
      RECT 108.411 108.166 110 110 ;
      RECT 108.273 108.304 110 110 ;
      RECT 108.365 108.212 110 110 ;
      RECT 108.319 108.258 110 110 ;
    LAYER MET3 SPACING 0.1 ;
      RECT -20 -20 3.325 110 ;
      RECT -20 -20 3.371 55.817 ;
      RECT -20 -20 3.417 55.771 ;
      RECT -20 -20 3.463 55.725 ;
      RECT -20 -20 3.509 55.679 ;
      RECT -20 -20 3.555 55.633 ;
      RECT -20 -20 3.601 55.587 ;
      RECT -20 -20 3.647 55.541 ;
      RECT -20 -20 3.693 55.495 ;
      RECT -20 -20 3.739 55.449 ;
      RECT -20 -20 3.785 55.403 ;
      RECT -20 -20 3.831 55.357 ;
      RECT -20 -20 3.877 55.311 ;
      RECT -20 -20 3.923 55.265 ;
      RECT -20 -20 3.969 55.219 ;
      RECT -20 -20 4.015 55.173 ;
      RECT -20 -20 4.061 55.127 ;
      RECT -20 -20 4.107 55.081 ;
      RECT -20 -20 4.153 55.035 ;
      RECT -20 -20 4.199 54.989 ;
      RECT -20 -20 4.245 54.943 ;
      RECT -20 -20 4.291 54.897 ;
      RECT -20 -20 4.337 54.851 ;
      RECT -20 -20 4.383 54.805 ;
      RECT -20 -20 4.429 54.759 ;
      RECT -20 -20 4.475 54.713 ;
      RECT -20 -20 4.521 54.667 ;
      RECT -20 -20 4.567 54.621 ;
      RECT -20 -20 4.613 54.575 ;
      RECT -20 -20 4.659 54.529 ;
      RECT -20 -20 4.705 54.483 ;
      RECT -20 -20 4.751 54.437 ;
      RECT -20 -20 4.797 54.391 ;
      RECT -20 -20 4.843 54.345 ;
      RECT -20 -20 4.889 54.299 ;
      RECT -20 -20 4.935 54.253 ;
      RECT -20 -20 4.981 54.207 ;
      RECT -20 -20 5.027 54.161 ;
      RECT -20 -20 5.073 54.115 ;
      RECT -20 -20 5.119 54.069 ;
      RECT -20 -20 5.165 54.023 ;
      RECT -20 -20 5.211 53.977 ;
      RECT -20 -20 5.257 53.931 ;
      RECT -20 -20 5.303 53.885 ;
      RECT -20 -20 5.349 53.839 ;
      RECT -20 -20 5.395 53.793 ;
      RECT -20 -20 5.441 53.747 ;
      RECT -20 -20 5.487 53.701 ;
      RECT -20 -20 5.533 53.655 ;
      RECT -20 -20 5.579 53.609 ;
      RECT -20 -20 5.625 53.563 ;
      RECT -20 -20 5.671 53.517 ;
      RECT -20 -20 5.717 53.471 ;
      RECT -20 -20 5.763 53.425 ;
      RECT -20 -20 5.809 53.379 ;
      RECT -20 -20 5.855 53.333 ;
      RECT -20 -20 5.901 53.287 ;
      RECT -20 -20 5.947 53.241 ;
      RECT -20 -20 5.993 53.195 ;
      RECT -20 -20 6.039 53.149 ;
      RECT -20 -20 6.085 53.103 ;
      RECT -20 -20 6.131 53.057 ;
      RECT -20 -20 6.177 53.011 ;
      RECT -20 -20 6.223 52.965 ;
      RECT -20 -20 6.269 52.919 ;
      RECT -20 -20 6.315 52.873 ;
      RECT -20 -20 6.361 52.827 ;
      RECT -20 -20 6.407 52.781 ;
      RECT -20 -20 6.453 52.735 ;
      RECT -20 -20 6.499 52.689 ;
      RECT -20 -20 6.545 52.643 ;
      RECT -20 -20 6.591 52.597 ;
      RECT -20 -20 6.637 52.551 ;
      RECT -20 -20 6.683 52.505 ;
      RECT -20 -20 6.729 52.459 ;
      RECT -20 -20 6.775 52.413 ;
      RECT -20 -20 6.821 52.367 ;
      RECT -20 -20 6.867 52.321 ;
      RECT -20 -20 6.913 52.275 ;
      RECT -20 -20 6.959 52.229 ;
      RECT -20 -20 7.005 52.183 ;
      RECT -20 -20 7.051 52.137 ;
      RECT -20 -20 7.097 52.091 ;
      RECT -20 -20 7.143 52.045 ;
      RECT -20 -20 7.189 51.999 ;
      RECT -20 -20 7.235 51.953 ;
      RECT -20 -20 7.281 51.907 ;
      RECT -20 -20 7.327 51.861 ;
      RECT -20 -20 7.373 51.815 ;
      RECT -20 -20 7.419 51.769 ;
      RECT -20 -20 7.465 51.723 ;
      RECT -20 -20 7.511 51.677 ;
      RECT -20 -20 7.557 51.631 ;
      RECT -20 -20 7.603 51.585 ;
      RECT -20 -20 7.649 51.539 ;
      RECT -20 -20 7.695 51.493 ;
      RECT -20 -20 7.741 51.447 ;
      RECT -20 -20 7.787 51.401 ;
      RECT -20 -20 7.833 51.355 ;
      RECT -20 -20 7.879 51.309 ;
      RECT -20 -20 7.925 51.263 ;
      RECT -20 -20 7.971 51.217 ;
      RECT -20 -20 8.017 51.171 ;
      RECT -20 -20 8.063 51.125 ;
      RECT -20 -20 8.109 51.079 ;
      RECT -20 -20 8.155 51.033 ;
      RECT -20 -20 8.201 50.987 ;
      RECT -20 -20 8.247 50.941 ;
      RECT -20 -20 8.293 50.895 ;
      RECT -20 -20 8.339 50.849 ;
      RECT -20 -20 8.385 50.803 ;
      RECT -20 -20 8.431 50.757 ;
      RECT -20 -20 8.477 50.711 ;
      RECT -20 -20 8.523 50.665 ;
      RECT -20 -20 8.569 50.619 ;
      RECT -20 -20 8.615 50.573 ;
      RECT -20 -20 8.661 50.527 ;
      RECT -20 -20 8.707 50.481 ;
      RECT -20 -20 8.753 50.435 ;
      RECT -20 -20 8.799 50.389 ;
      RECT -20 -20 8.845 50.343 ;
      RECT -20 -20 8.891 50.297 ;
      RECT -20 -20 8.937 50.251 ;
      RECT -20 -20 8.983 50.205 ;
      RECT -20 -20 9.029 50.159 ;
      RECT -20 -20 9.075 50.113 ;
      RECT -20 -20 9.121 50.067 ;
      RECT -20 -20 9.167 50.021 ;
      RECT -20 -20 9.213 49.975 ;
      RECT -20 -20 9.259 49.929 ;
      RECT -20 -20 9.305 49.883 ;
      RECT -20 -20 9.351 49.837 ;
      RECT -20 -20 9.397 49.791 ;
      RECT -20 -20 9.443 49.745 ;
      RECT -20 -20 9.489 49.699 ;
      RECT -20 -20 9.535 49.653 ;
      RECT -20 -20 9.581 49.607 ;
      RECT -20 -20 9.627 49.561 ;
      RECT -20 -20 9.673 49.515 ;
      RECT -20 -20 9.719 49.469 ;
      RECT -20 -20 9.765 49.423 ;
      RECT -20 -20 9.811 49.377 ;
      RECT -20 -20 9.857 49.331 ;
      RECT -20 -20 9.903 49.285 ;
      RECT -20 -20 9.949 49.239 ;
      RECT -20 -20 9.995 49.193 ;
      RECT -20 -20 10.041 49.147 ;
      RECT -20 -20 10.087 49.101 ;
      RECT -20 -20 10.133 49.055 ;
      RECT -20 -20 10.179 49.009 ;
      RECT -20 -20 10.225 48.963 ;
      RECT -20 -20 10.271 48.917 ;
      RECT -20 -20 10.317 48.871 ;
      RECT -20 -20 10.363 48.825 ;
      RECT -20 -20 10.409 48.779 ;
      RECT -20 -20 10.455 48.733 ;
      RECT -20 -20 10.501 48.687 ;
      RECT -20 -20 10.547 48.641 ;
      RECT -20 -20 10.593 48.595 ;
      RECT -20 -20 10.639 48.549 ;
      RECT -20 -20 10.685 48.503 ;
      RECT -20 -20 10.731 48.457 ;
      RECT -20 -20 10.777 48.411 ;
      RECT -20 -20 10.823 48.365 ;
      RECT -20 -20 10.869 48.319 ;
      RECT -20 -20 10.915 48.273 ;
      RECT -20 -20 10.961 48.227 ;
      RECT -20 -20 11.007 48.181 ;
      RECT -20 -20 11.053 48.135 ;
      RECT -20 -20 11.099 48.089 ;
      RECT -20 -20 11.145 48.043 ;
      RECT -20 -20 11.191 47.997 ;
      RECT -20 -20 11.237 47.951 ;
      RECT -20 -20 11.283 47.905 ;
      RECT -20 -20 11.329 47.859 ;
      RECT -20 -20 11.375 47.813 ;
      RECT -20 -20 11.421 47.767 ;
      RECT -20 -20 11.467 47.721 ;
      RECT -20 -20 11.513 47.675 ;
      RECT -20 -20 11.559 47.629 ;
      RECT -20 -20 11.605 47.583 ;
      RECT -20 -20 11.651 47.537 ;
      RECT -20 -20 11.697 47.491 ;
      RECT -20 -20 11.743 47.445 ;
      RECT -20 -20 11.789 47.399 ;
      RECT -20 -20 11.835 47.353 ;
      RECT -20 -20 11.881 47.307 ;
      RECT -20 -20 11.927 47.261 ;
      RECT -20 -20 11.973 47.215 ;
      RECT -20 -20 12.019 47.169 ;
      RECT -20 -20 12.065 47.123 ;
      RECT -20 -20 12.111 47.077 ;
      RECT -20 -20 12.157 47.031 ;
      RECT -20 -20 12.203 46.985 ;
      RECT -20 -20 12.249 46.939 ;
      RECT -20 -20 12.295 46.893 ;
      RECT -20 -20 12.341 46.847 ;
      RECT -20 -20 12.387 46.801 ;
      RECT -20 -20 12.433 46.755 ;
      RECT -20 -20 12.479 46.709 ;
      RECT -20 -20 12.525 46.663 ;
      RECT -20 -20 12.571 46.617 ;
      RECT -20 -20 12.617 46.571 ;
      RECT -20 -20 12.663 46.525 ;
      RECT -20 -20 12.709 46.479 ;
      RECT -20 -20 12.755 46.433 ;
      RECT -20 -20 12.801 46.387 ;
      RECT -20 -20 12.847 46.341 ;
      RECT -20 -20 12.893 46.295 ;
      RECT -20 -20 12.939 46.249 ;
      RECT -20 -20 12.985 46.203 ;
      RECT -20 -20 13.031 46.157 ;
      RECT -20 -20 13.077 46.111 ;
      RECT -20 -20 13.123 46.065 ;
      RECT -20 -20 13.169 46.019 ;
      RECT -20 -20 13.215 45.973 ;
      RECT -20 -20 13.261 45.927 ;
      RECT -20 -20 13.307 45.881 ;
      RECT -20 -20 13.353 45.835 ;
      RECT -20 -20 13.399 45.789 ;
      RECT -20 -20 13.445 45.743 ;
      RECT -20 -20 13.491 45.697 ;
      RECT -20 -20 13.537 45.651 ;
      RECT -20 -20 13.583 45.605 ;
      RECT -20 -20 13.629 45.559 ;
      RECT -20 -20 13.675 45.513 ;
      RECT -20 -20 13.721 45.467 ;
      RECT -20 -20 13.767 45.421 ;
      RECT -20 -20 13.813 45.375 ;
      RECT -20 -20 13.859 45.329 ;
      RECT -20 -20 13.905 45.283 ;
      RECT -20 -20 13.951 45.237 ;
      RECT -20 -20 13.997 45.191 ;
      RECT -20 -20 14.043 45.145 ;
      RECT -20 -20 14.089 45.099 ;
      RECT -20 -20 14.135 45.053 ;
      RECT -20 -20 14.181 45.007 ;
      RECT -20 -20 14.227 44.961 ;
      RECT -20 -20 14.273 44.915 ;
      RECT -20 -20 14.319 44.869 ;
      RECT -20 -20 14.365 44.823 ;
      RECT -20 -20 14.411 44.777 ;
      RECT -20 -20 14.457 44.731 ;
      RECT -20 -20 14.503 44.685 ;
      RECT -20 -20 14.549 44.639 ;
      RECT -20 -20 14.595 44.593 ;
      RECT -20 -20 14.641 44.547 ;
      RECT -20 -20 14.687 44.501 ;
      RECT -20 -20 14.733 44.455 ;
      RECT -20 -20 14.779 44.409 ;
      RECT -20 -20 14.825 44.363 ;
      RECT -20 -20 14.871 44.317 ;
      RECT -20 -20 14.917 44.271 ;
      RECT -20 -20 14.963 44.225 ;
      RECT -20 -20 15.009 44.179 ;
      RECT -20 -20 15.055 44.133 ;
      RECT -20 -20 15.101 44.087 ;
      RECT -20 -20 15.147 44.041 ;
      RECT -20 -20 15.193 43.995 ;
      RECT -20 -20 15.239 43.949 ;
      RECT -20 -20 15.285 43.903 ;
      RECT -20 -20 15.325 43.86 ;
      RECT -20 -20 15.371 43.817 ;
      RECT -20 -20 15.417 43.771 ;
      RECT -20 -20 15.463 43.725 ;
      RECT -20 -20 15.509 43.679 ;
      RECT -20 -20 15.555 43.633 ;
      RECT -20 -20 15.601 43.587 ;
      RECT -20 -20 15.647 43.541 ;
      RECT -20 -20 15.693 43.495 ;
      RECT -20 -20 15.739 43.449 ;
      RECT -20 -20 15.785 43.403 ;
      RECT -20 -20 15.831 43.357 ;
      RECT -20 -20 15.877 43.311 ;
      RECT -20 -20 15.923 43.265 ;
      RECT -20 -20 15.969 43.219 ;
      RECT -20 -20 16.015 43.173 ;
      RECT -20 -20 16.061 43.127 ;
      RECT -20 -20 16.107 43.081 ;
      RECT -20 -20 16.153 43.035 ;
      RECT -20 -20 16.199 42.989 ;
      RECT -20 -20 16.245 42.943 ;
      RECT -20 -20 16.291 42.897 ;
      RECT -20 -20 16.337 42.851 ;
      RECT -20 -20 16.383 42.805 ;
      RECT -20 -20 16.429 42.759 ;
      RECT -20 -20 16.475 42.713 ;
      RECT -20 -20 16.521 42.667 ;
      RECT -20 -20 16.567 42.621 ;
      RECT -20 -20 16.613 42.575 ;
      RECT -20 -20 16.659 42.529 ;
      RECT -20 -20 16.705 42.483 ;
      RECT -20 -20 16.751 42.437 ;
      RECT -20 -20 16.797 42.391 ;
      RECT -20 -20 16.843 42.345 ;
      RECT -20 -20 16.889 42.299 ;
      RECT -20 -20 16.935 42.253 ;
      RECT -20 -20 16.981 42.207 ;
      RECT -20 -20 17.027 42.161 ;
      RECT -20 -20 17.073 42.115 ;
      RECT -20 -20 17.119 42.069 ;
      RECT -20 -20 17.165 42.023 ;
      RECT -20 -20 17.211 41.977 ;
      RECT -20 -20 17.257 41.931 ;
      RECT -20 -20 17.303 41.885 ;
      RECT -20 -20 17.349 41.839 ;
      RECT -20 -20 17.395 41.793 ;
      RECT -20 -20 17.441 41.747 ;
      RECT -20 -20 17.487 41.701 ;
      RECT -20 -20 17.533 41.655 ;
      RECT -20 -20 17.579 41.609 ;
      RECT -20 -20 17.625 41.563 ;
      RECT -20 -20 17.671 41.517 ;
      RECT -20 -20 17.717 41.471 ;
      RECT -20 -20 17.763 41.425 ;
      RECT -20 -20 17.809 41.379 ;
      RECT -20 -20 17.855 41.333 ;
      RECT -20 -20 17.901 41.287 ;
      RECT -20 -20 17.947 41.241 ;
      RECT -20 -20 17.993 41.195 ;
      RECT -20 -20 18.039 41.149 ;
      RECT -20 -20 18.085 41.103 ;
      RECT -20 -20 18.131 41.057 ;
      RECT -20 -20 18.177 41.011 ;
      RECT -20 -20 18.223 40.965 ;
      RECT -20 -20 18.269 40.919 ;
      RECT -20 -20 18.315 40.873 ;
      RECT -20 -20 18.361 40.827 ;
      RECT -20 -20 18.407 40.781 ;
      RECT -20 -20 18.453 40.735 ;
      RECT -20 -20 18.499 40.689 ;
      RECT -20 -20 18.545 40.643 ;
      RECT -20 -20 18.591 40.597 ;
      RECT -20 -20 18.637 40.551 ;
      RECT -20 -20 18.683 40.505 ;
      RECT -20 -20 18.729 40.459 ;
      RECT -20 -20 18.775 40.413 ;
      RECT -20 -20 18.821 40.367 ;
      RECT -20 -20 18.867 40.321 ;
      RECT -20 -20 18.913 40.275 ;
      RECT -20 -20 18.959 40.229 ;
      RECT -20 -20 19.005 40.183 ;
      RECT -20 -20 19.051 40.137 ;
      RECT -20 -20 19.097 40.091 ;
      RECT -20 -20 19.143 40.045 ;
      RECT -20 -20 19.189 39.999 ;
      RECT -20 -20 19.235 39.953 ;
      RECT -20 -20 19.281 39.907 ;
      RECT -20 -20 19.327 39.861 ;
      RECT -20 -20 19.373 39.815 ;
      RECT -20 -20 19.419 39.769 ;
      RECT -20 -20 19.465 39.723 ;
      RECT -20 -20 19.511 39.677 ;
      RECT -20 -20 19.557 39.631 ;
      RECT -20 -20 19.603 39.585 ;
      RECT -20 -20 19.649 39.539 ;
      RECT -20 -20 19.695 39.493 ;
      RECT -20 -20 19.741 39.447 ;
      RECT -20 -20 19.787 39.401 ;
      RECT -20 -20 19.833 39.355 ;
      RECT -20 -20 19.879 39.309 ;
      RECT -20 -20 19.925 39.263 ;
      RECT -20 -20 19.971 39.217 ;
      RECT -20 -20 20.017 39.171 ;
      RECT -20 -20 20.063 39.125 ;
      RECT -20 -20 20.109 39.079 ;
      RECT -20 -20 20.155 39.033 ;
      RECT -20 -20 20.201 38.987 ;
      RECT -20 -20 20.247 38.941 ;
      RECT -20 -20 20.293 38.895 ;
      RECT -20 -20 20.339 38.849 ;
      RECT -20 -20 20.385 38.803 ;
      RECT -20 -20 20.431 38.757 ;
      RECT -20 -20 20.477 38.711 ;
      RECT -20 -20 20.523 38.665 ;
      RECT -20 -20 20.569 38.619 ;
      RECT -20 -20 20.615 38.573 ;
      RECT -20 -20 20.661 38.527 ;
      RECT -20 -20 20.707 38.481 ;
      RECT -20 -20 20.753 38.435 ;
      RECT -20 -20 20.799 38.389 ;
      RECT -20 -20 20.845 38.343 ;
      RECT -20 -20 20.891 38.297 ;
      RECT -20 -20 20.937 38.251 ;
      RECT -20 -20 20.983 38.205 ;
      RECT -20 -20 21.029 38.159 ;
      RECT -20 -20 21.075 38.113 ;
      RECT -20 -20 21.121 38.067 ;
      RECT -20 -20 21.167 38.021 ;
      RECT -20 -20 21.213 37.975 ;
      RECT -20 -20 21.259 37.929 ;
      RECT -20 -20 21.305 37.883 ;
      RECT -20 -20 21.351 37.837 ;
      RECT -20 -20 21.397 37.791 ;
      RECT -20 -20 21.443 37.745 ;
      RECT -20 -20 21.489 37.699 ;
      RECT -20 -20 21.535 37.653 ;
      RECT -20 -20 21.581 37.607 ;
      RECT -20 -20 21.627 37.561 ;
      RECT -20 -20 21.673 37.515 ;
      RECT -20 -20 21.719 37.469 ;
      RECT -20 -20 21.765 37.423 ;
      RECT -20 -20 21.811 37.377 ;
      RECT -20 -20 21.857 37.331 ;
      RECT -20 -20 21.903 37.285 ;
      RECT -20 -20 21.949 37.239 ;
      RECT -20 -20 21.995 37.193 ;
      RECT -20 -20 22.041 37.147 ;
      RECT -20 -20 22.087 37.101 ;
      RECT -20 -20 22.133 37.055 ;
      RECT -20 -20 22.179 37.009 ;
      RECT -20 -20 22.225 36.963 ;
      RECT -20 -20 22.271 36.917 ;
      RECT -20 -20 22.317 36.871 ;
      RECT -20 -20 22.363 36.825 ;
      RECT -20 -20 22.409 36.779 ;
      RECT -20 -20 22.455 36.733 ;
      RECT -20 -20 22.501 36.687 ;
      RECT -20 -20 22.547 36.641 ;
      RECT -20 -20 22.593 36.595 ;
      RECT -20 -20 22.639 36.549 ;
      RECT -20 -20 22.685 36.503 ;
      RECT -20 -20 22.731 36.457 ;
      RECT -20 -20 22.777 36.411 ;
      RECT -20 -20 22.823 36.365 ;
      RECT -20 -20 22.869 36.319 ;
      RECT -20 -20 22.915 36.273 ;
      RECT -20 -20 22.961 36.227 ;
      RECT -20 -20 23.007 36.181 ;
      RECT -20 -20 23.053 36.135 ;
      RECT -20 -20 23.099 36.089 ;
      RECT -20 -20 23.145 36.043 ;
      RECT -20 -20 23.191 35.997 ;
      RECT -20 -20 23.237 35.951 ;
      RECT -20 -20 23.283 35.905 ;
      RECT -20 -20 23.329 35.859 ;
      RECT -20 -20 23.375 35.813 ;
      RECT -20 -20 23.421 35.767 ;
      RECT -20 -20 23.467 35.721 ;
      RECT -20 -20 23.513 35.675 ;
      RECT -20 -20 23.559 35.629 ;
      RECT -20 -20 23.605 35.583 ;
      RECT -20 -20 23.651 35.537 ;
      RECT -20 -20 23.697 35.491 ;
      RECT -20 -20 23.743 35.445 ;
      RECT -20 -20 23.789 35.399 ;
      RECT -20 -20 23.835 35.353 ;
      RECT -20 -20 23.881 35.307 ;
      RECT -20 -20 23.927 35.261 ;
      RECT -20 -20 23.973 35.215 ;
      RECT -20 -20 24.019 35.169 ;
      RECT -20 -20 24.065 35.123 ;
      RECT -20 -20 24.111 35.077 ;
      RECT -20 -20 24.157 35.031 ;
      RECT -20 -20 24.203 34.985 ;
      RECT -20 -20 24.249 34.939 ;
      RECT -20 -20 24.295 34.893 ;
      RECT -20 -20 24.341 34.847 ;
      RECT -20 -20 24.387 34.801 ;
      RECT -20 -20 24.433 34.755 ;
      RECT -20 -20 24.479 34.709 ;
      RECT -20 -20 24.525 34.663 ;
      RECT -20 -20 24.571 34.617 ;
      RECT -20 -20 24.617 34.571 ;
      RECT -20 -20 24.663 34.525 ;
      RECT -20 -20 24.709 34.479 ;
      RECT -20 -20 24.755 34.433 ;
      RECT -20 -20 24.801 34.387 ;
      RECT -20 -20 24.847 34.341 ;
      RECT -20 -20 24.893 34.295 ;
      RECT -20 -20 24.939 34.249 ;
      RECT -20 -20 24.985 34.203 ;
      RECT -20 -20 25.031 34.157 ;
      RECT -20 -20 25.077 34.111 ;
      RECT -20 -20 25.123 34.065 ;
      RECT -20 -20 25.169 34.019 ;
      RECT -20 -20 25.215 33.973 ;
      RECT -20 -20 25.261 33.927 ;
      RECT -20 -20 25.307 33.881 ;
      RECT -20 -20 25.353 33.835 ;
      RECT -20 -20 25.399 33.789 ;
      RECT -20 -20 25.445 33.743 ;
      RECT -20 -20 25.491 33.697 ;
      RECT -20 -20 25.537 33.651 ;
      RECT -20 -20 25.583 33.605 ;
      RECT -20 -20 25.629 33.559 ;
      RECT -20 -20 25.675 33.513 ;
      RECT -20 -20 25.721 33.467 ;
      RECT -20 -20 25.767 33.421 ;
      RECT -20 -20 25.813 33.375 ;
      RECT -20 -20 25.859 33.329 ;
      RECT -20 -20 25.905 33.283 ;
      RECT -20 -20 25.951 33.237 ;
      RECT -20 -20 25.997 33.191 ;
      RECT -20 -20 26.043 33.145 ;
      RECT -20 -20 26.089 33.099 ;
      RECT -20 -20 26.135 33.053 ;
      RECT -20 -20 26.181 33.007 ;
      RECT -20 -20 26.227 32.961 ;
      RECT -20 -20 26.273 32.915 ;
      RECT -20 -20 26.319 32.869 ;
      RECT -20 -20 26.365 32.823 ;
      RECT -20 -20 26.411 32.777 ;
      RECT -20 -20 26.457 32.731 ;
      RECT -20 -20 26.503 32.685 ;
      RECT -20 -20 26.549 32.639 ;
      RECT -20 -20 26.595 32.593 ;
      RECT -20 -20 26.641 32.547 ;
      RECT -20 -20 26.687 32.501 ;
      RECT -20 -20 26.733 32.455 ;
      RECT -20 -20 26.779 32.409 ;
      RECT -20 -20 26.825 32.363 ;
      RECT -20 -20 26.871 32.317 ;
      RECT -20 -20 26.917 32.271 ;
      RECT -20 -20 26.963 32.225 ;
      RECT -20 -20 27.009 32.179 ;
      RECT -20 -20 27.055 32.133 ;
      RECT -20 -20 27.101 32.087 ;
      RECT -20 -20 27.147 32.041 ;
      RECT -20 -20 27.193 31.995 ;
      RECT -20 -20 27.239 31.949 ;
      RECT -20 -20 27.285 31.903 ;
      RECT -20 -20 27.331 31.857 ;
      RECT -20 -20 27.377 31.811 ;
      RECT -20 -20 27.423 31.765 ;
      RECT -20 -20 27.469 31.719 ;
      RECT -20 -20 27.515 31.673 ;
      RECT -20 -20 27.561 31.627 ;
      RECT -20 -20 27.607 31.581 ;
      RECT -20 -20 27.653 31.535 ;
      RECT -20 -20 27.699 31.489 ;
      RECT -20 -20 27.745 31.443 ;
      RECT -20 -20 27.791 31.397 ;
      RECT -20 -20 27.837 31.351 ;
      RECT -20 -20 27.883 31.305 ;
      RECT -20 -20 27.929 31.259 ;
      RECT -20 -20 27.975 31.213 ;
      RECT -20 -20 28.021 31.167 ;
      RECT -20 -20 28.067 31.121 ;
      RECT -20 -20 28.113 31.075 ;
      RECT -20 -20 28.159 31.029 ;
      RECT -20 -20 28.205 30.983 ;
      RECT -20 -20 28.251 30.937 ;
      RECT -20 -20 28.297 30.891 ;
      RECT -20 -20 28.343 30.845 ;
      RECT -20 -20 28.389 30.799 ;
      RECT -20 -20 28.435 30.753 ;
      RECT -20 -20 28.481 30.707 ;
      RECT -20 -20 28.527 30.661 ;
      RECT -20 -20 28.573 30.615 ;
      RECT -20 -20 28.619 30.569 ;
      RECT -20 -20 28.665 30.523 ;
      RECT -20 -20 28.711 30.477 ;
      RECT -20 -20 28.757 30.431 ;
      RECT -20 -20 28.803 30.385 ;
      RECT -20 -20 28.849 30.339 ;
      RECT -20 -20 28.895 30.293 ;
      RECT -20 -20 28.941 30.247 ;
      RECT -20 -20 28.987 30.201 ;
      RECT -20 -20 29.033 30.155 ;
      RECT -20 -20 29.079 30.109 ;
      RECT -20 -20 29.125 30.063 ;
      RECT -20 -20 29.171 30.017 ;
      RECT -20 -20 29.217 29.971 ;
      RECT -20 -20 29.263 29.925 ;
      RECT -20 -20 29.309 29.879 ;
      RECT -20 -20 29.355 29.833 ;
      RECT -20 -20 29.401 29.787 ;
      RECT -20 -20 29.447 29.741 ;
      RECT -20 -20 29.493 29.695 ;
      RECT -20 -20 29.539 29.649 ;
      RECT -20 -20 29.585 29.603 ;
      RECT -20 -20 29.631 29.557 ;
      RECT -20 -20 29.677 29.511 ;
      RECT -20 -20 29.723 29.465 ;
      RECT -20 -20 29.769 29.419 ;
      RECT -20 -20 29.815 29.373 ;
      RECT -20 -20 29.861 29.327 ;
      RECT -20 -20 29.907 29.281 ;
      RECT -20 -20 29.953 29.235 ;
      RECT -20 -20 29.999 29.189 ;
      RECT -20 -20 30.045 29.143 ;
      RECT -20 -20 30.091 29.097 ;
      RECT -20 -20 30.137 29.051 ;
      RECT -20 -20 30.183 29.005 ;
      RECT -20 -20 30.229 28.959 ;
      RECT -20 -20 30.275 28.913 ;
      RECT -20 -20 30.321 28.867 ;
      RECT -20 -20 30.367 28.821 ;
      RECT -20 -20 30.413 28.775 ;
      RECT -20 -20 30.459 28.729 ;
      RECT -20 -20 30.505 28.683 ;
      RECT -20 -20 30.551 28.637 ;
      RECT -20 -20 30.597 28.591 ;
      RECT -20 -20 30.643 28.545 ;
      RECT -20 -20 30.689 28.499 ;
      RECT -20 -20 30.735 28.453 ;
      RECT -20 -20 30.781 28.407 ;
      RECT -20 -20 30.827 28.361 ;
      RECT -20 -20 30.873 28.315 ;
      RECT -20 -20 30.919 28.269 ;
      RECT -20 -20 30.965 28.223 ;
      RECT -20 -20 31.011 28.177 ;
      RECT -20 -20 31.057 28.131 ;
      RECT -20 -20 31.103 28.085 ;
      RECT -20 -20 31.149 28.039 ;
      RECT -20 -20 31.195 27.993 ;
      RECT -20 -20 31.241 27.947 ;
      RECT -20 -20 31.287 27.901 ;
      RECT -20 -20 31.333 27.855 ;
      RECT -20 -20 31.379 27.809 ;
      RECT -20 -20 31.425 27.763 ;
      RECT -20 -20 31.471 27.717 ;
      RECT -20 -20 31.517 27.671 ;
      RECT -20 -20 31.563 27.625 ;
      RECT -20 -20 31.609 27.579 ;
      RECT -20 -20 31.655 27.533 ;
      RECT -20 -20 31.701 27.487 ;
      RECT -20 -20 31.747 27.441 ;
      RECT -20 -20 31.793 27.395 ;
      RECT -20 -20 31.839 27.349 ;
      RECT -20 -20 31.885 27.303 ;
      RECT -20 -20 31.931 27.257 ;
      RECT -20 -20 31.977 27.211 ;
      RECT -20 -20 32.023 27.165 ;
      RECT -20 -20 32.069 27.119 ;
      RECT -20 -20 32.115 27.073 ;
      RECT -20 -20 32.161 27.027 ;
      RECT -20 -20 32.207 26.981 ;
      RECT -20 -20 32.253 26.935 ;
      RECT -20 -20 32.299 26.889 ;
      RECT -20 -20 32.345 26.843 ;
      RECT -20 -20 32.391 26.797 ;
      RECT -20 -20 32.437 26.751 ;
      RECT -20 -20 32.483 26.705 ;
      RECT -20 -20 32.529 26.659 ;
      RECT -20 -20 32.575 26.613 ;
      RECT -20 -20 32.621 26.567 ;
      RECT -20 -20 32.667 26.521 ;
      RECT -20 -20 32.713 26.475 ;
      RECT -20 -20 32.759 26.429 ;
      RECT -20 -20 32.805 26.383 ;
      RECT -20 -20 32.851 26.337 ;
      RECT -20 -20 32.897 26.291 ;
      RECT -20 -20 32.943 26.245 ;
      RECT -20 -20 32.989 26.199 ;
      RECT -20 -20 33.035 26.153 ;
      RECT -20 -20 33.081 26.107 ;
      RECT -20 -20 33.127 26.061 ;
      RECT -20 -20 33.173 26.015 ;
      RECT -20 -20 33.219 25.969 ;
      RECT -20 -20 33.265 25.923 ;
      RECT -20 -20 33.311 25.877 ;
      RECT -20 -20 33.357 25.831 ;
      RECT -20 -20 33.403 25.785 ;
      RECT -20 -20 33.449 25.739 ;
      RECT -20 -20 33.495 25.693 ;
      RECT -20 -20 33.541 25.647 ;
      RECT -20 -20 33.587 25.601 ;
      RECT -20 -20 33.633 25.555 ;
      RECT -20 -20 33.679 25.509 ;
      RECT -20 -20 33.725 25.463 ;
      RECT -20 -20 33.771 25.417 ;
      RECT -20 -20 33.817 25.371 ;
      RECT -20 -20 33.863 25.325 ;
      RECT -20 -20 33.909 25.279 ;
      RECT -20 -20 33.955 25.233 ;
      RECT -20 -20 34.001 25.187 ;
      RECT -20 -20 34.047 25.141 ;
      RECT -20 -20 34.093 25.095 ;
      RECT -20 -20 34.139 25.049 ;
      RECT -20 -20 34.185 25.003 ;
      RECT -20 -20 34.231 24.957 ;
      RECT -20 -20 34.277 24.911 ;
      RECT -20 -20 34.323 24.865 ;
      RECT -20 -20 34.369 24.819 ;
      RECT -20 -20 34.415 24.773 ;
      RECT -20 -20 34.461 24.727 ;
      RECT -20 -20 34.507 24.681 ;
      RECT -20 -20 34.553 24.635 ;
      RECT -20 -20 34.599 24.589 ;
      RECT -20 -20 34.645 24.543 ;
      RECT -20 -20 34.691 24.497 ;
      RECT -20 -20 34.737 24.451 ;
      RECT -20 -20 34.783 24.405 ;
      RECT -20 -20 34.829 24.359 ;
      RECT -20 -20 34.875 24.313 ;
      RECT -20 -20 34.921 24.267 ;
      RECT -20 -20 34.967 24.221 ;
      RECT -20 -20 35.013 24.175 ;
      RECT -20 -20 35.059 24.129 ;
      RECT -20 -20 35.105 24.083 ;
      RECT -20 -20 35.151 24.037 ;
      RECT -20 -20 35.197 23.991 ;
      RECT -20 -20 35.243 23.945 ;
      RECT -20 -20 35.289 23.899 ;
      RECT -20 -20 35.335 23.853 ;
      RECT -20 -20 35.381 23.807 ;
      RECT -20 -20 35.427 23.761 ;
      RECT -20 -20 35.473 23.715 ;
      RECT -20 -20 35.519 23.669 ;
      RECT -20 -20 35.565 23.623 ;
      RECT -20 -20 35.611 23.577 ;
      RECT -20 -20 35.657 23.531 ;
      RECT -20 -20 35.703 23.485 ;
      RECT -20 -20 35.749 23.439 ;
      RECT -20 -20 35.795 23.393 ;
      RECT -20 -20 35.841 23.347 ;
      RECT -20 -20 35.887 23.301 ;
      RECT -20 -20 35.933 23.255 ;
      RECT -20 -20 35.979 23.209 ;
      RECT -20 -20 36.025 23.163 ;
      RECT -20 -20 36.071 23.117 ;
      RECT -20 -20 36.117 23.071 ;
      RECT -20 -20 36.163 23.025 ;
      RECT -20 -20 36.209 22.979 ;
      RECT -20 -20 36.255 22.933 ;
      RECT -20 -20 36.301 22.887 ;
      RECT -20 -20 36.347 22.841 ;
      RECT -20 -20 36.393 22.795 ;
      RECT -20 -20 36.439 22.749 ;
      RECT -20 -20 36.485 22.703 ;
      RECT -20 -20 36.531 22.657 ;
      RECT -20 -20 36.577 22.611 ;
      RECT -20 -20 36.623 22.565 ;
      RECT -20 -20 36.669 22.519 ;
      RECT -20 -20 36.715 22.473 ;
      RECT -20 -20 36.761 22.427 ;
      RECT -20 -20 36.807 22.381 ;
      RECT -20 -20 36.853 22.335 ;
      RECT -20 -20 36.899 22.289 ;
      RECT -20 -20 36.945 22.243 ;
      RECT -20 -20 36.991 22.197 ;
      RECT -20 -20 37.037 22.151 ;
      RECT -20 -20 37.083 22.105 ;
      RECT -20 -20 37.129 22.059 ;
      RECT -20 -20 37.175 22.013 ;
      RECT -20 -20 37.221 21.967 ;
      RECT -20 -20 37.267 21.921 ;
      RECT -20 -20 37.313 21.875 ;
      RECT -20 -20 37.359 21.829 ;
      RECT -20 -20 37.405 21.783 ;
      RECT -20 -20 37.451 21.737 ;
      RECT -20 -20 37.497 21.691 ;
      RECT -20 -20 37.543 21.645 ;
      RECT -20 -20 37.589 21.599 ;
      RECT -20 -20 37.635 21.553 ;
      RECT -20 -20 37.681 21.507 ;
      RECT -20 -20 37.727 21.461 ;
      RECT -20 -20 37.773 21.415 ;
      RECT -20 -20 37.819 21.369 ;
      RECT -20 -20 37.865 21.323 ;
      RECT -20 -20 37.911 21.277 ;
      RECT -20 -20 37.957 21.231 ;
      RECT -20 -20 38.003 21.185 ;
      RECT -20 -20 38.049 21.139 ;
      RECT -20 -20 38.095 21.093 ;
      RECT -20 -20 38.141 21.047 ;
      RECT -20 -20 38.187 21.001 ;
      RECT -20 -20 38.233 20.955 ;
      RECT -20 -20 38.279 20.909 ;
      RECT -20 -20 38.325 20.863 ;
      RECT -20 -20 38.371 20.817 ;
      RECT -20 -20 38.417 20.771 ;
      RECT -20 -20 38.463 20.725 ;
      RECT -20 -20 38.509 20.679 ;
      RECT -20 -20 38.555 20.633 ;
      RECT -20 -20 38.601 20.587 ;
      RECT -20 -20 38.647 20.541 ;
      RECT -20 -20 38.693 20.495 ;
      RECT -20 -20 38.739 20.449 ;
      RECT -20 -20 38.785 20.403 ;
      RECT -20 -20 38.831 20.357 ;
      RECT -20 -20 38.877 20.311 ;
      RECT -20 -20 38.923 20.265 ;
      RECT -20 -20 38.969 20.219 ;
      RECT -20 -20 39.015 20.173 ;
      RECT -20 -20 39.061 20.127 ;
      RECT -20 -20 39.107 20.081 ;
      RECT -20 -20 39.153 20.035 ;
      RECT -20 -20 39.199 19.989 ;
      RECT -20 -20 39.245 19.943 ;
      RECT -20 -20 39.291 19.897 ;
      RECT -20 -20 39.337 19.851 ;
      RECT -20 -20 39.383 19.805 ;
      RECT -20 -20 39.429 19.759 ;
      RECT -20 -20 39.475 19.713 ;
      RECT -20 -20 39.521 19.667 ;
      RECT -20 -20 39.567 19.621 ;
      RECT -20 -20 39.613 19.575 ;
      RECT -20 -20 39.659 19.529 ;
      RECT -20 -20 39.705 19.483 ;
      RECT -20 -20 39.751 19.437 ;
      RECT -20 -20 39.797 19.391 ;
      RECT -20 -20 39.843 19.345 ;
      RECT -20 -20 39.889 19.299 ;
      RECT -20 -20 39.935 19.253 ;
      RECT -20 -20 39.981 19.207 ;
      RECT -20 -20 40.027 19.161 ;
      RECT -20 -20 40.073 19.115 ;
      RECT -20 -20 40.119 19.069 ;
      RECT -20 -20 40.165 19.023 ;
      RECT -20 -20 40.211 18.977 ;
      RECT -20 -20 40.257 18.931 ;
      RECT -20 -20 40.303 18.885 ;
      RECT -20 -20 40.349 18.839 ;
      RECT -20 -20 40.395 18.793 ;
      RECT -20 -20 40.441 18.747 ;
      RECT -20 -20 40.487 18.701 ;
      RECT -20 -20 40.533 18.655 ;
      RECT -20 -20 40.579 18.609 ;
      RECT -20 -20 40.625 18.563 ;
      RECT -20 -20 40.671 18.517 ;
      RECT -20 -20 40.717 18.471 ;
      RECT -20 -20 40.763 18.425 ;
      RECT -20 -20 40.809 18.379 ;
      RECT -20 -20 40.855 18.333 ;
      RECT -20 -20 40.901 18.287 ;
      RECT -20 -20 40.947 18.241 ;
      RECT -20 -20 40.993 18.195 ;
      RECT -20 -20 41.039 18.149 ;
      RECT -20 -20 41.085 18.103 ;
      RECT -20 -20 41.131 18.057 ;
      RECT -20 -20 41.177 18.011 ;
      RECT -20 -20 41.223 17.965 ;
      RECT -20 -20 41.269 17.919 ;
      RECT -20 -20 41.315 17.873 ;
      RECT -20 -20 41.361 17.827 ;
      RECT -20 -20 41.407 17.781 ;
      RECT -20 -20 41.453 17.735 ;
      RECT -20 -20 41.499 17.689 ;
      RECT -20 -20 41.545 17.643 ;
      RECT -20 -20 41.591 17.597 ;
      RECT -20 -20 41.637 17.551 ;
      RECT -20 -20 41.683 17.505 ;
      RECT -20 -20 41.729 17.459 ;
      RECT -20 -20 41.775 17.413 ;
      RECT -20 -20 41.821 17.367 ;
      RECT -20 -20 41.867 17.321 ;
      RECT -20 -20 41.913 17.275 ;
      RECT -20 -20 41.959 17.229 ;
      RECT -20 -20 42.005 17.183 ;
      RECT -20 -20 42.051 17.137 ;
      RECT -20 -20 42.097 17.091 ;
      RECT -20 -20 42.143 17.045 ;
      RECT -20 -20 42.189 16.999 ;
      RECT -20 -20 42.235 16.953 ;
      RECT -20 -20 42.281 16.907 ;
      RECT -20 -20 42.327 16.861 ;
      RECT -20 -20 42.373 16.815 ;
      RECT -20 -20 42.419 16.769 ;
      RECT -20 -20 42.465 16.723 ;
      RECT -20 -20 42.511 16.677 ;
      RECT -20 -20 42.557 16.631 ;
      RECT -20 -20 42.603 16.585 ;
      RECT -20 -20 42.649 16.539 ;
      RECT -20 -20 42.695 16.493 ;
      RECT -20 -20 42.741 16.447 ;
      RECT -20 -20 42.787 16.401 ;
      RECT -20 -20 42.833 16.355 ;
      RECT -20 -20 42.879 16.309 ;
      RECT -20 -20 42.925 16.263 ;
      RECT -20 -20 42.971 16.217 ;
      RECT -20 -20 43.017 16.171 ;
      RECT -20 -20 43.063 16.125 ;
      RECT -20 -20 43.109 16.079 ;
      RECT -20 -20 43.155 16.033 ;
      RECT -20 -20 43.201 15.987 ;
      RECT -20 -20 43.247 15.941 ;
      RECT -20 -20 43.293 15.895 ;
      RECT -20 -20 43.339 15.849 ;
      RECT -20 -20 43.385 15.803 ;
      RECT -20 -20 43.431 15.757 ;
      RECT -20 -20 43.477 15.711 ;
      RECT -20 -20 43.523 15.665 ;
      RECT -20 -20 43.569 15.619 ;
      RECT -20 -20 43.615 15.573 ;
      RECT -20 -20 43.661 15.527 ;
      RECT -20 -20 43.707 15.481 ;
      RECT -20 -20 43.753 15.435 ;
      RECT -20 -20 43.799 15.389 ;
      RECT -20 -20 43.845 15.343 ;
      RECT -20 -20 43.891 15.297 ;
      RECT -20 -20 43.937 15.251 ;
      RECT -20 -20 43.983 15.205 ;
      RECT -20 -20 44.029 15.159 ;
      RECT -20 -20 44.075 15.113 ;
      RECT -20 -20 44.121 15.067 ;
      RECT -20 -20 44.167 15.021 ;
      RECT -20 -20 44.213 14.975 ;
      RECT -20 -20 44.259 14.929 ;
      RECT -20 -20 44.305 14.883 ;
      RECT -20 -20 44.351 14.837 ;
      RECT -20 -20 44.397 14.791 ;
      RECT -20 -20 44.443 14.745 ;
      RECT -20 -20 44.489 14.699 ;
      RECT -20 -20 44.535 14.653 ;
      RECT -20 -20 44.581 14.607 ;
      RECT -20 -20 44.627 14.561 ;
      RECT -20 -20 44.673 14.515 ;
      RECT -20 -20 44.719 14.469 ;
      RECT -20 -20 44.765 14.423 ;
      RECT -20 -20 44.811 14.377 ;
      RECT -20 -20 44.857 14.331 ;
      RECT -20 -20 44.903 14.285 ;
      RECT -20 -20 44.949 14.239 ;
      RECT -20 -20 44.995 14.193 ;
      RECT -20 -20 45.041 14.147 ;
      RECT -20 -20 45.087 14.101 ;
      RECT -20 -20 45.133 14.055 ;
      RECT -20 -20 45.179 14.009 ;
      RECT -20 -20 45.225 13.963 ;
      RECT -20 -20 45.271 13.917 ;
      RECT -20 -20 45.317 13.871 ;
      RECT -20 -20 45.363 13.825 ;
      RECT -20 -20 45.409 13.779 ;
      RECT -20 -20 45.455 13.733 ;
      RECT -20 -20 45.501 13.687 ;
      RECT -20 -20 45.547 13.641 ;
      RECT -20 -20 45.593 13.595 ;
      RECT -20 -20 45.639 13.549 ;
      RECT -20 -20 45.685 13.503 ;
      RECT -20 -20 45.731 13.457 ;
      RECT -20 -20 45.777 13.411 ;
      RECT -20 -20 45.823 13.365 ;
      RECT -20 -20 45.869 13.319 ;
      RECT -20 -20 45.915 13.273 ;
      RECT -20 -20 45.961 13.227 ;
      RECT -20 -20 46.007 13.181 ;
      RECT -20 -20 46.053 13.135 ;
      RECT -20 -20 46.099 13.089 ;
      RECT -20 -20 46.145 13.043 ;
      RECT -20 -20 46.191 12.997 ;
      RECT -20 -20 46.237 12.951 ;
      RECT -20 -20 46.283 12.905 ;
      RECT -20 -20 46.329 12.859 ;
      RECT -20 -20 46.375 12.813 ;
      RECT -20 -20 46.421 12.767 ;
      RECT -20 -20 46.467 12.721 ;
      RECT -20 -20 46.513 12.675 ;
      RECT -20 -20 46.559 12.629 ;
      RECT -20 -20 46.605 12.583 ;
      RECT -20 -20 46.651 12.537 ;
      RECT -20 -20 46.697 12.491 ;
      RECT -20 -20 46.743 12.445 ;
      RECT -20 -20 46.789 12.399 ;
      RECT -20 -20 46.835 12.353 ;
      RECT -20 -20 46.881 12.307 ;
      RECT -20 -20 46.927 12.261 ;
      RECT -20 -20 46.973 12.215 ;
      RECT -20 -20 47.019 12.169 ;
      RECT -20 -20 47.065 12.123 ;
      RECT -20 -20 47.111 12.077 ;
      RECT -20 -20 47.157 12.031 ;
      RECT -20 -20 47.203 11.985 ;
      RECT -20 -20 47.249 11.939 ;
      RECT -20 -20 47.295 11.893 ;
      RECT -20 -20 47.341 11.847 ;
      RECT -20 -20 47.387 11.801 ;
      RECT -20 -20 47.433 11.755 ;
      RECT -20 -20 47.479 11.709 ;
      RECT -20 -20 47.525 11.663 ;
      RECT -20 -20 47.571 11.617 ;
      RECT -20 -20 47.617 11.571 ;
      RECT -20 -20 47.663 11.525 ;
      RECT -20 -20 47.709 11.479 ;
      RECT -20 -20 47.755 11.433 ;
      RECT -20 -20 47.801 11.387 ;
      RECT -20 -20 47.847 11.341 ;
      RECT -20 -20 47.893 11.295 ;
      RECT -20 -20 47.939 11.249 ;
      RECT -20 -20 47.985 11.203 ;
      RECT -20 -20 48.031 11.157 ;
      RECT -20 -20 48.077 11.111 ;
      RECT -20 -20 48.123 11.065 ;
      RECT -20 -20 48.169 11.019 ;
      RECT -20 -20 48.215 10.973 ;
      RECT -20 -20 48.261 10.927 ;
      RECT -20 -20 48.307 10.881 ;
      RECT -20 -20 48.353 10.835 ;
      RECT -20 -20 48.399 10.789 ;
      RECT -20 -20 48.445 10.743 ;
      RECT -20 -20 48.491 10.697 ;
      RECT -20 -20 48.537 10.651 ;
      RECT -20 -20 48.583 10.605 ;
      RECT -20 -20 48.629 10.559 ;
      RECT -20 -20 48.675 10.513 ;
      RECT -20 -20 48.721 10.467 ;
      RECT -20 -20 48.767 10.421 ;
      RECT -20 -20 48.813 10.375 ;
      RECT -20 -20 48.859 10.329 ;
      RECT -20 -20 48.905 10.283 ;
      RECT -20 -20 48.951 10.237 ;
      RECT -20 -20 48.997 10.191 ;
      RECT -20 -20 49.043 10.145 ;
      RECT -20 -20 49.089 10.099 ;
      RECT -20 -20 49.135 10.053 ;
      RECT -20 -20 49.181 10.007 ;
      RECT -20 -20 49.227 9.961 ;
      RECT -20 -20 49.273 9.915 ;
      RECT -20 -20 49.319 9.869 ;
      RECT -20 -20 49.365 9.823 ;
      RECT -20 -20 49.411 9.777 ;
      RECT -20 -20 49.457 9.731 ;
      RECT -20 -20 49.503 9.685 ;
      RECT -20 -20 49.549 9.639 ;
      RECT -20 -20 49.595 9.593 ;
      RECT -20 -20 49.641 9.547 ;
      RECT -20 -20 49.687 9.501 ;
      RECT -20 -20 49.733 9.455 ;
      RECT -20 -20 49.779 9.409 ;
      RECT -20 -20 49.825 9.363 ;
      RECT -20 -20 49.871 9.317 ;
      RECT -20 -20 49.917 9.271 ;
      RECT -20 -20 49.963 9.225 ;
      RECT -20 -20 50.009 9.179 ;
      RECT -20 -20 50.055 9.133 ;
      RECT -20 -20 50.101 9.087 ;
      RECT -20 -20 50.147 9.041 ;
      RECT -20 -20 50.193 8.995 ;
      RECT -20 -20 50.239 8.949 ;
      RECT -20 -20 50.285 8.903 ;
      RECT -20 -20 50.331 8.857 ;
      RECT -20 -20 50.377 8.811 ;
      RECT -20 -20 50.423 8.765 ;
      RECT -20 -20 50.469 8.719 ;
      RECT -20 -20 50.515 8.673 ;
      RECT -20 -20 50.561 8.627 ;
      RECT -20 -20 50.607 8.581 ;
      RECT -20 -20 50.653 8.535 ;
      RECT -20 -20 50.699 8.489 ;
      RECT -20 -20 50.745 8.443 ;
      RECT -20 -20 50.791 8.397 ;
      RECT -20 -20 50.837 8.351 ;
      RECT -20 -20 50.883 8.305 ;
      RECT -20 -20 50.929 8.259 ;
      RECT -20 -20 50.975 8.213 ;
      RECT -20 -20 51.021 8.167 ;
      RECT -20 -20 51.067 8.121 ;
      RECT -20 -20 51.113 8.075 ;
      RECT -20 -20 51.159 8.029 ;
      RECT -20 -20 51.205 7.983 ;
      RECT -20 -20 51.251 7.937 ;
      RECT -20 -20 51.297 7.891 ;
      RECT -20 -20 51.343 7.845 ;
      RECT -20 -20 51.389 7.799 ;
      RECT -20 -20 51.435 7.753 ;
      RECT -20 -20 51.481 7.707 ;
      RECT -20 -20 51.527 7.661 ;
      RECT -20 -20 51.573 7.615 ;
      RECT -20 -20 51.619 7.569 ;
      RECT -20 -20 51.665 7.523 ;
      RECT -20 -20 51.711 7.477 ;
      RECT -20 -20 51.757 7.431 ;
      RECT -20 -20 51.803 7.385 ;
      RECT -20 -20 51.849 7.339 ;
      RECT -20 -20 51.895 7.293 ;
      RECT -20 -20 51.941 7.247 ;
      RECT -20 -20 51.987 7.201 ;
      RECT -20 -20 52.033 7.155 ;
      RECT -20 -20 52.079 7.109 ;
      RECT -20 -20 52.125 7.063 ;
      RECT -20 -20 52.171 7.017 ;
      RECT -20 -20 52.217 6.971 ;
      RECT -20 -20 52.263 6.925 ;
      RECT -20 -20 52.309 6.879 ;
      RECT -20 -20 52.355 6.833 ;
      RECT -20 -20 52.401 6.787 ;
      RECT -20 -20 52.447 6.741 ;
      RECT -20 -20 52.493 6.695 ;
      RECT -20 -20 52.539 6.649 ;
      RECT -20 -20 52.585 6.603 ;
      RECT -20 -20 52.631 6.557 ;
      RECT -20 -20 52.677 6.511 ;
      RECT -20 -20 52.723 6.465 ;
      RECT -20 -20 52.769 6.419 ;
      RECT -20 -20 52.815 6.373 ;
      RECT -20 -20 52.861 6.327 ;
      RECT -20 -20 52.907 6.281 ;
      RECT -20 -20 52.953 6.235 ;
      RECT -20 -20 52.999 6.189 ;
      RECT -20 -20 53.045 6.143 ;
      RECT -20 -20 53.091 6.097 ;
      RECT -20 -20 53.137 6.051 ;
      RECT -20 -20 53.183 6.005 ;
      RECT -20 -20 53.229 5.959 ;
      RECT -20 -20 53.275 5.913 ;
      RECT -20 -20 53.321 5.867 ;
      RECT -20 -20 53.367 5.821 ;
      RECT -20 -20 53.413 5.775 ;
      RECT -20 -20 53.459 5.729 ;
      RECT -20 -20 53.505 5.683 ;
      RECT -20 -20 53.551 5.637 ;
      RECT -20 -20 53.597 5.591 ;
      RECT -20 -20 53.643 5.545 ;
      RECT -20 -20 53.689 5.499 ;
      RECT -20 -20 53.735 5.453 ;
      RECT -20 -20 53.781 5.407 ;
      RECT -20 -20 53.827 5.361 ;
      RECT -20 -20 53.873 5.315 ;
      RECT -20 -20 53.919 5.269 ;
      RECT -20 -20 53.965 5.223 ;
      RECT -20 -20 54.011 5.177 ;
      RECT -20 -20 54.057 5.131 ;
      RECT -20 -20 54.103 5.085 ;
      RECT -20 -20 54.149 5.039 ;
      RECT -20 -20 54.195 4.993 ;
      RECT -20 -20 54.241 4.947 ;
      RECT -20 -20 54.287 4.901 ;
      RECT -20 -20 54.333 4.855 ;
      RECT -20 -20 54.379 4.809 ;
      RECT -20 -20 54.425 4.763 ;
      RECT -20 -20 54.471 4.717 ;
      RECT -20 -20 54.517 4.671 ;
      RECT -20 -20 54.563 4.625 ;
      RECT -20 -20 54.609 4.579 ;
      RECT -20 -20 54.655 4.533 ;
      RECT -20 -20 54.701 4.487 ;
      RECT -20 -20 54.747 4.441 ;
      RECT -20 -20 54.793 4.395 ;
      RECT -20 -20 54.839 4.349 ;
      RECT -20 -20 54.885 4.303 ;
      RECT -20 -20 54.931 4.257 ;
      RECT -20 -20 54.977 4.211 ;
      RECT -20 -20 55.023 4.165 ;
      RECT -20 -20 55.069 4.119 ;
      RECT -20 -20 55.115 4.073 ;
      RECT -20 -20 55.161 4.027 ;
      RECT -20 -20 55.207 3.981 ;
      RECT -20 -20 55.253 3.935 ;
      RECT -20 -20 55.299 3.889 ;
      RECT -20 -20 55.345 3.843 ;
      RECT -20 -20 55.391 3.797 ;
      RECT -20 -20 55.437 3.751 ;
      RECT -20 -20 55.483 3.705 ;
      RECT -20 -20 55.529 3.659 ;
      RECT -20 -20 55.575 3.613 ;
      RECT -20 -20 55.621 3.567 ;
      RECT -20 -20 55.667 3.521 ;
      RECT -20 -20 55.713 3.475 ;
      RECT -20 -20 55.759 3.429 ;
      RECT -20 -20 55.805 3.383 ;
      RECT -20 -20 55.84 3.342 ;
      RECT -20 -20 110 3.325 ;
      RECT 15.675 61.137 16.825 110 ;
      RECT 15.675 61.137 16.871 62.567 ;
      RECT 15.675 61.137 16.917 62.521 ;
      RECT 15.675 61.137 16.963 62.475 ;
      RECT 15.675 61.137 17.009 62.429 ;
      RECT 15.675 61.137 17.055 62.383 ;
      RECT 15.675 61.137 17.101 62.337 ;
      RECT 15.675 61.137 17.147 62.291 ;
      RECT 15.675 61.137 17.193 62.245 ;
      RECT 15.675 61.137 17.239 62.199 ;
      RECT 15.675 61.137 17.285 62.153 ;
      RECT 15.675 61.137 17.331 62.107 ;
      RECT 15.675 61.137 17.377 62.061 ;
      RECT 15.675 61.137 17.423 62.015 ;
      RECT 15.675 61.137 17.469 61.969 ;
      RECT 15.675 61.137 17.515 61.923 ;
      RECT 15.675 61.137 17.561 61.877 ;
      RECT 15.675 61.137 17.607 61.831 ;
      RECT 15.675 61.137 17.653 61.785 ;
      RECT 15.675 61.137 17.699 61.739 ;
      RECT 15.675 61.137 17.745 61.693 ;
      RECT 15.675 61.137 17.791 61.647 ;
      RECT 15.675 61.137 17.837 61.601 ;
      RECT 15.675 61.137 17.883 61.555 ;
      RECT 15.675 61.137 17.929 61.509 ;
      RECT 15.675 61.137 17.975 61.463 ;
      RECT 15.675 61.137 18.021 61.417 ;
      RECT 15.675 61.137 18.067 61.371 ;
      RECT 15.675 61.137 18.113 61.325 ;
      RECT 15.675 61.137 18.159 61.279 ;
      RECT 15.675 61.137 18.205 61.233 ;
      RECT 15.675 61.137 18.251 61.187 ;
      RECT 15.721 61.091 18.297 61.141 ;
      RECT 15.767 61.045 18.343 61.095 ;
      RECT 15.813 60.999 18.389 61.049 ;
      RECT 15.859 60.953 18.435 61.003 ;
      RECT 15.905 60.907 18.481 60.957 ;
      RECT 15.951 60.861 18.527 60.911 ;
      RECT 15.997 60.815 18.573 60.865 ;
      RECT 16.043 60.769 18.619 60.819 ;
      RECT 16.089 60.723 18.665 60.773 ;
      RECT 16.135 60.677 18.711 60.727 ;
      RECT 16.181 60.631 18.757 60.681 ;
      RECT 16.227 60.585 18.803 60.635 ;
      RECT 16.273 60.539 18.849 60.589 ;
      RECT 16.319 60.493 18.895 60.543 ;
      RECT 16.365 60.447 18.941 60.497 ;
      RECT 16.411 60.401 18.987 60.451 ;
      RECT 16.457 60.355 19.033 60.405 ;
      RECT 16.503 60.309 19.079 60.359 ;
      RECT 16.549 60.263 19.125 60.313 ;
      RECT 16.595 60.217 19.171 60.267 ;
      RECT 16.641 60.171 19.217 60.221 ;
      RECT 16.687 60.125 19.263 60.175 ;
      RECT 16.733 60.079 19.309 60.129 ;
      RECT 16.779 60.033 19.355 60.083 ;
      RECT 16.825 59.987 19.401 60.037 ;
      RECT 16.871 59.941 19.447 59.991 ;
      RECT 16.917 59.895 19.493 59.945 ;
      RECT 16.963 59.849 19.539 59.899 ;
      RECT 17.009 59.803 19.585 59.853 ;
      RECT 17.055 59.757 19.631 59.807 ;
      RECT 17.101 59.711 19.677 59.761 ;
      RECT 17.147 59.665 19.723 59.715 ;
      RECT 17.193 59.619 19.769 59.669 ;
      RECT 17.239 59.573 19.815 59.623 ;
      RECT 17.285 59.527 19.861 59.577 ;
      RECT 17.331 59.481 19.907 59.531 ;
      RECT 17.377 59.435 19.953 59.485 ;
      RECT 17.423 59.389 19.999 59.439 ;
      RECT 17.469 59.343 20.045 59.393 ;
      RECT 17.515 59.297 20.091 59.347 ;
      RECT 17.561 59.251 20.137 59.301 ;
      RECT 17.607 59.205 20.183 59.255 ;
      RECT 17.653 59.159 20.229 59.209 ;
      RECT 17.699 59.113 20.275 59.163 ;
      RECT 17.745 59.067 20.321 59.117 ;
      RECT 17.791 59.021 20.367 59.071 ;
      RECT 17.837 58.975 20.413 59.025 ;
      RECT 17.883 58.929 20.459 58.979 ;
      RECT 17.929 58.883 20.505 58.933 ;
      RECT 17.975 58.837 20.551 58.887 ;
      RECT 18.021 58.791 20.597 58.841 ;
      RECT 18.067 58.745 20.643 58.795 ;
      RECT 18.113 58.699 20.689 58.749 ;
      RECT 18.159 58.653 20.735 58.703 ;
      RECT 18.205 58.607 20.781 58.657 ;
      RECT 18.251 58.561 20.827 58.611 ;
      RECT 18.297 58.515 20.873 58.565 ;
      RECT 18.343 58.469 20.919 58.519 ;
      RECT 18.389 58.423 20.965 58.473 ;
      RECT 18.435 58.377 21.011 58.427 ;
      RECT 18.481 58.331 21.057 58.381 ;
      RECT 18.527 58.285 21.103 58.335 ;
      RECT 18.573 58.239 21.149 58.289 ;
      RECT 18.619 58.193 21.195 58.243 ;
      RECT 18.665 58.147 21.241 58.197 ;
      RECT 18.711 58.101 21.287 58.151 ;
      RECT 18.757 58.055 21.333 58.105 ;
      RECT 18.803 58.009 21.379 58.059 ;
      RECT 18.849 57.963 21.425 58.013 ;
      RECT 18.895 57.917 21.471 57.967 ;
      RECT 18.941 57.871 21.517 57.921 ;
      RECT 18.987 57.825 21.563 57.875 ;
      RECT 19.033 57.779 21.609 57.829 ;
      RECT 19.079 57.733 21.655 57.783 ;
      RECT 19.125 57.687 21.701 57.737 ;
      RECT 19.171 57.641 21.747 57.691 ;
      RECT 19.217 57.595 21.793 57.645 ;
      RECT 19.263 57.549 21.839 57.599 ;
      RECT 19.309 57.503 21.885 57.553 ;
      RECT 19.355 57.457 21.931 57.507 ;
      RECT 19.401 57.411 21.977 57.461 ;
      RECT 19.447 57.365 22.023 57.415 ;
      RECT 19.493 57.319 22.069 57.369 ;
      RECT 19.539 57.273 22.115 57.323 ;
      RECT 19.585 57.227 22.161 57.277 ;
      RECT 19.631 57.181 22.207 57.231 ;
      RECT 19.677 57.135 22.253 57.185 ;
      RECT 19.723 57.089 22.299 57.139 ;
      RECT 19.769 57.043 22.345 57.093 ;
      RECT 19.815 56.997 22.391 57.047 ;
      RECT 19.861 56.951 22.437 57.001 ;
      RECT 19.907 56.905 22.483 56.955 ;
      RECT 19.953 56.859 22.529 56.909 ;
      RECT 19.999 56.813 22.575 56.863 ;
      RECT 20.045 56.767 22.621 56.817 ;
      RECT 20.091 56.721 22.667 56.771 ;
      RECT 20.137 56.675 22.713 56.725 ;
      RECT 20.183 56.629 22.759 56.679 ;
      RECT 20.229 56.583 22.805 56.633 ;
      RECT 20.275 56.537 22.851 56.587 ;
      RECT 20.321 56.491 22.897 56.541 ;
      RECT 20.367 56.445 22.943 56.495 ;
      RECT 20.413 56.399 22.989 56.449 ;
      RECT 20.459 56.353 23.035 56.403 ;
      RECT 20.505 56.307 23.081 56.357 ;
      RECT 20.551 56.261 23.127 56.311 ;
      RECT 20.597 56.215 23.173 56.265 ;
      RECT 20.643 56.169 23.219 56.219 ;
      RECT 20.689 56.123 23.265 56.173 ;
      RECT 20.735 56.077 23.311 56.127 ;
      RECT 20.781 56.031 23.357 56.081 ;
      RECT 20.827 55.985 23.403 56.035 ;
      RECT 20.873 55.939 23.449 55.989 ;
      RECT 20.919 55.893 23.495 55.943 ;
      RECT 20.965 55.847 23.541 55.897 ;
      RECT 21.011 55.801 23.587 55.851 ;
      RECT 21.057 55.755 23.633 55.805 ;
      RECT 21.103 55.709 23.679 55.759 ;
      RECT 21.149 55.663 23.725 55.713 ;
      RECT 21.195 55.617 23.771 55.667 ;
      RECT 21.241 55.571 23.817 55.621 ;
      RECT 21.287 55.525 23.863 55.575 ;
      RECT 21.333 55.479 23.909 55.529 ;
      RECT 21.379 55.433 23.955 55.483 ;
      RECT 21.425 55.387 24.001 55.437 ;
      RECT 21.471 55.341 24.047 55.391 ;
      RECT 21.517 55.295 24.093 55.345 ;
      RECT 21.563 55.249 24.139 55.299 ;
      RECT 21.609 55.203 24.185 55.253 ;
      RECT 21.655 55.157 24.231 55.207 ;
      RECT 21.701 55.111 24.277 55.161 ;
      RECT 21.747 55.065 24.323 55.115 ;
      RECT 21.793 55.019 24.369 55.069 ;
      RECT 21.839 54.973 24.415 55.023 ;
      RECT 21.885 54.927 24.461 54.977 ;
      RECT 21.931 54.881 24.507 54.931 ;
      RECT 21.977 54.835 24.553 54.885 ;
      RECT 22.023 54.789 24.599 54.839 ;
      RECT 22.069 54.743 24.645 54.793 ;
      RECT 22.115 54.697 24.691 54.747 ;
      RECT 22.161 54.651 24.737 54.701 ;
      RECT 22.207 54.605 24.783 54.655 ;
      RECT 22.253 54.559 24.829 54.609 ;
      RECT 22.299 54.513 24.875 54.563 ;
      RECT 22.345 54.467 24.921 54.517 ;
      RECT 22.391 54.421 24.967 54.471 ;
      RECT 22.437 54.375 25.013 54.425 ;
      RECT 22.483 54.329 25.059 54.379 ;
      RECT 22.529 54.283 25.105 54.333 ;
      RECT 22.575 54.237 25.151 54.287 ;
      RECT 22.621 54.191 25.197 54.241 ;
      RECT 22.667 54.145 25.243 54.195 ;
      RECT 22.713 54.099 25.289 54.149 ;
      RECT 22.759 54.053 25.335 54.103 ;
      RECT 22.805 54.007 25.381 54.057 ;
      RECT 22.851 53.961 25.427 54.011 ;
      RECT 22.897 53.915 25.473 53.965 ;
      RECT 22.943 53.869 25.519 53.919 ;
      RECT 22.989 53.823 25.565 53.873 ;
      RECT 23.035 53.777 25.611 53.827 ;
      RECT 23.081 53.731 25.657 53.781 ;
      RECT 23.127 53.685 25.703 53.735 ;
      RECT 23.173 53.639 25.749 53.689 ;
      RECT 23.219 53.593 25.795 53.643 ;
      RECT 23.265 53.547 25.841 53.597 ;
      RECT 23.311 53.501 25.887 53.551 ;
      RECT 23.357 53.455 25.933 53.505 ;
      RECT 23.403 53.409 25.979 53.459 ;
      RECT 23.449 53.363 26.025 53.413 ;
      RECT 23.495 53.317 26.071 53.367 ;
      RECT 23.541 53.271 26.117 53.321 ;
      RECT 23.587 53.225 26.163 53.275 ;
      RECT 23.633 53.179 26.209 53.229 ;
      RECT 23.679 53.133 26.255 53.183 ;
      RECT 23.725 53.087 26.301 53.137 ;
      RECT 23.771 53.041 26.347 53.091 ;
      RECT 23.817 52.995 26.393 53.045 ;
      RECT 23.863 52.949 26.439 52.999 ;
      RECT 23.909 52.903 26.485 52.953 ;
      RECT 23.955 52.857 26.531 52.907 ;
      RECT 24.001 52.811 26.577 52.861 ;
      RECT 24.047 52.765 26.623 52.815 ;
      RECT 24.093 52.719 26.669 52.769 ;
      RECT 24.139 52.673 26.715 52.723 ;
      RECT 24.185 52.627 26.761 52.677 ;
      RECT 24.231 52.581 26.807 52.631 ;
      RECT 24.277 52.535 26.853 52.585 ;
      RECT 24.323 52.489 26.899 52.539 ;
      RECT 24.369 52.443 26.945 52.493 ;
      RECT 24.415 52.397 26.991 52.447 ;
      RECT 24.461 52.351 27.037 52.401 ;
      RECT 24.507 52.305 27.083 52.355 ;
      RECT 24.553 52.259 27.129 52.309 ;
      RECT 24.599 52.213 27.175 52.263 ;
      RECT 24.645 52.167 27.221 52.217 ;
      RECT 24.691 52.121 27.267 52.171 ;
      RECT 24.737 52.075 27.313 52.125 ;
      RECT 24.783 52.029 27.359 52.079 ;
      RECT 24.829 51.983 27.405 52.033 ;
      RECT 24.875 51.937 27.451 51.987 ;
      RECT 24.921 51.891 27.497 51.941 ;
      RECT 24.967 51.845 27.543 51.895 ;
      RECT 25.013 51.799 27.589 51.849 ;
      RECT 25.059 51.753 27.635 51.803 ;
      RECT 25.105 51.707 27.681 51.757 ;
      RECT 25.151 51.661 27.727 51.711 ;
      RECT 25.197 51.615 27.773 51.665 ;
      RECT 25.243 51.569 27.819 51.619 ;
      RECT 25.289 51.523 27.865 51.573 ;
      RECT 25.335 51.477 27.911 51.527 ;
      RECT 25.381 51.431 27.957 51.481 ;
      RECT 25.427 51.385 28.003 51.435 ;
      RECT 25.473 51.339 28.049 51.389 ;
      RECT 25.519 51.293 28.095 51.343 ;
      RECT 25.565 51.247 28.141 51.297 ;
      RECT 25.611 51.201 28.187 51.251 ;
      RECT 25.657 51.155 28.233 51.205 ;
      RECT 25.703 51.109 28.279 51.159 ;
      RECT 25.749 51.063 28.325 51.113 ;
      RECT 25.795 51.017 28.371 51.067 ;
      RECT 25.841 50.971 28.417 51.021 ;
      RECT 25.887 50.925 28.463 50.975 ;
      RECT 25.933 50.879 28.509 50.929 ;
      RECT 25.979 50.833 28.555 50.883 ;
      RECT 26.025 50.787 28.601 50.837 ;
      RECT 26.071 50.741 28.647 50.791 ;
      RECT 26.117 50.695 28.693 50.745 ;
      RECT 26.163 50.649 28.739 50.699 ;
      RECT 26.209 50.603 28.785 50.653 ;
      RECT 26.255 50.557 28.825 50.61 ;
      RECT 26.301 50.511 28.871 50.567 ;
      RECT 26.347 50.465 28.917 50.521 ;
      RECT 26.393 50.419 28.963 50.475 ;
      RECT 26.439 50.373 29.009 50.429 ;
      RECT 26.485 50.327 29.055 50.383 ;
      RECT 26.531 50.281 29.101 50.337 ;
      RECT 26.577 50.235 29.147 50.291 ;
      RECT 26.623 50.189 29.193 50.245 ;
      RECT 26.669 50.143 29.239 50.199 ;
      RECT 26.715 50.097 29.285 50.153 ;
      RECT 26.761 50.051 29.331 50.107 ;
      RECT 26.807 50.005 29.377 50.061 ;
      RECT 26.853 49.959 29.423 50.015 ;
      RECT 26.899 49.913 29.469 49.969 ;
      RECT 26.945 49.867 29.515 49.923 ;
      RECT 26.991 49.821 29.561 49.877 ;
      RECT 27.037 49.775 29.607 49.831 ;
      RECT 27.083 49.729 29.653 49.785 ;
      RECT 27.129 49.683 29.699 49.739 ;
      RECT 27.175 49.637 29.745 49.693 ;
      RECT 27.221 49.591 29.791 49.647 ;
      RECT 27.267 49.545 29.837 49.601 ;
      RECT 27.313 49.499 29.883 49.555 ;
      RECT 27.359 49.453 29.929 49.509 ;
      RECT 27.405 49.407 29.975 49.463 ;
      RECT 27.451 49.361 30.021 49.417 ;
      RECT 27.497 49.315 30.067 49.371 ;
      RECT 27.543 49.269 30.113 49.325 ;
      RECT 27.589 49.223 30.159 49.279 ;
      RECT 27.635 49.177 30.205 49.233 ;
      RECT 27.681 49.131 30.251 49.187 ;
      RECT 27.727 49.085 30.297 49.141 ;
      RECT 27.773 49.039 30.343 49.095 ;
      RECT 27.819 48.993 30.389 49.049 ;
      RECT 27.865 48.947 30.435 49.003 ;
      RECT 27.911 48.901 30.481 48.957 ;
      RECT 27.957 48.855 30.527 48.911 ;
      RECT 28.003 48.809 30.573 48.865 ;
      RECT 28.049 48.763 30.619 48.819 ;
      RECT 28.095 48.717 30.665 48.773 ;
      RECT 28.141 48.671 30.711 48.727 ;
      RECT 28.187 48.625 30.757 48.681 ;
      RECT 28.233 48.579 30.803 48.635 ;
      RECT 28.279 48.533 30.849 48.589 ;
      RECT 28.325 48.487 30.895 48.543 ;
      RECT 28.371 48.441 30.941 48.497 ;
      RECT 28.417 48.395 30.987 48.451 ;
      RECT 28.463 48.349 31.033 48.405 ;
      RECT 28.509 48.303 31.079 48.359 ;
      RECT 28.555 48.257 31.125 48.313 ;
      RECT 28.601 48.211 31.171 48.267 ;
      RECT 28.647 48.165 31.217 48.221 ;
      RECT 28.693 48.119 31.263 48.175 ;
      RECT 28.739 48.073 31.309 48.129 ;
      RECT 28.785 48.027 31.355 48.083 ;
      RECT 28.831 47.981 31.401 48.037 ;
      RECT 28.877 47.935 31.447 47.991 ;
      RECT 28.923 47.889 31.493 47.945 ;
      RECT 28.969 47.843 31.539 47.899 ;
      RECT 29.015 47.797 31.585 47.853 ;
      RECT 29.061 47.751 31.631 47.807 ;
      RECT 29.107 47.705 31.677 47.761 ;
      RECT 29.153 47.659 31.723 47.715 ;
      RECT 29.199 47.613 31.769 47.669 ;
      RECT 29.245 47.567 31.815 47.623 ;
      RECT 29.291 47.521 31.861 47.577 ;
      RECT 29.337 47.475 31.907 47.531 ;
      RECT 29.383 47.429 31.953 47.485 ;
      RECT 29.429 47.383 31.999 47.439 ;
      RECT 29.475 47.337 32.045 47.393 ;
      RECT 29.521 47.291 32.091 47.347 ;
      RECT 29.567 47.245 32.137 47.301 ;
      RECT 29.613 47.199 32.183 47.255 ;
      RECT 29.659 47.153 32.229 47.209 ;
      RECT 29.705 47.107 32.275 47.163 ;
      RECT 29.751 47.061 32.321 47.117 ;
      RECT 29.797 47.015 32.367 47.071 ;
      RECT 29.843 46.969 32.413 47.025 ;
      RECT 29.889 46.923 32.459 46.979 ;
      RECT 29.935 46.877 32.505 46.933 ;
      RECT 29.981 46.831 32.551 46.887 ;
      RECT 30.027 46.785 32.597 46.841 ;
      RECT 30.073 46.739 32.643 46.795 ;
      RECT 30.119 46.693 32.689 46.749 ;
      RECT 30.165 46.647 32.735 46.703 ;
      RECT 30.211 46.601 32.781 46.657 ;
      RECT 30.257 46.555 32.827 46.611 ;
      RECT 30.303 46.509 32.873 46.565 ;
      RECT 30.349 46.463 32.919 46.519 ;
      RECT 30.395 46.417 32.965 46.473 ;
      RECT 30.441 46.371 33.011 46.427 ;
      RECT 30.487 46.325 33.057 46.381 ;
      RECT 30.533 46.279 33.103 46.335 ;
      RECT 30.579 46.233 33.149 46.289 ;
      RECT 30.625 46.187 33.195 46.243 ;
      RECT 30.671 46.141 33.241 46.197 ;
      RECT 30.717 46.095 33.287 46.151 ;
      RECT 30.763 46.049 33.333 46.105 ;
      RECT 30.809 46.003 33.379 46.059 ;
      RECT 30.855 45.957 33.425 46.013 ;
      RECT 30.901 45.911 33.471 45.967 ;
      RECT 30.947 45.865 33.517 45.921 ;
      RECT 30.993 45.819 33.563 45.875 ;
      RECT 31.039 45.773 33.609 45.829 ;
      RECT 31.085 45.727 33.655 45.783 ;
      RECT 31.131 45.681 33.701 45.737 ;
      RECT 31.177 45.635 33.747 45.691 ;
      RECT 31.223 45.589 33.793 45.645 ;
      RECT 31.269 45.543 33.839 45.599 ;
      RECT 31.315 45.497 33.885 45.553 ;
      RECT 31.361 45.451 33.931 45.507 ;
      RECT 31.407 45.405 33.977 45.461 ;
      RECT 31.453 45.359 34.023 45.415 ;
      RECT 31.499 45.313 34.069 45.369 ;
      RECT 31.545 45.267 34.115 45.323 ;
      RECT 31.591 45.221 34.161 45.277 ;
      RECT 31.637 45.175 34.207 45.231 ;
      RECT 31.683 45.129 34.253 45.185 ;
      RECT 31.729 45.083 34.299 45.139 ;
      RECT 31.775 45.037 34.345 45.093 ;
      RECT 31.821 44.991 34.391 45.047 ;
      RECT 31.867 44.945 34.437 45.001 ;
      RECT 31.913 44.899 34.483 44.955 ;
      RECT 31.959 44.853 34.529 44.909 ;
      RECT 32.005 44.807 34.575 44.863 ;
      RECT 32.051 44.761 34.621 44.817 ;
      RECT 32.097 44.715 34.667 44.771 ;
      RECT 32.143 44.669 34.713 44.725 ;
      RECT 32.189 44.623 34.759 44.679 ;
      RECT 32.235 44.577 34.805 44.633 ;
      RECT 32.281 44.531 34.851 44.587 ;
      RECT 32.327 44.485 34.897 44.541 ;
      RECT 32.373 44.439 34.943 44.495 ;
      RECT 32.419 44.393 34.989 44.449 ;
      RECT 32.465 44.347 35.035 44.403 ;
      RECT 32.511 44.301 35.081 44.357 ;
      RECT 32.557 44.255 35.127 44.311 ;
      RECT 32.603 44.209 35.173 44.265 ;
      RECT 32.649 44.163 35.219 44.219 ;
      RECT 32.695 44.117 35.265 44.173 ;
      RECT 32.741 44.071 35.311 44.127 ;
      RECT 32.787 44.025 35.357 44.081 ;
      RECT 32.833 43.979 35.403 44.035 ;
      RECT 32.879 43.933 35.449 43.989 ;
      RECT 32.925 43.887 35.495 43.943 ;
      RECT 32.971 43.841 35.541 43.897 ;
      RECT 33.017 43.795 35.587 43.851 ;
      RECT 33.063 43.749 35.633 43.805 ;
      RECT 33.109 43.703 35.679 43.759 ;
      RECT 33.155 43.657 35.725 43.713 ;
      RECT 33.201 43.611 35.771 43.667 ;
      RECT 33.247 43.565 35.817 43.621 ;
      RECT 33.293 43.519 35.863 43.575 ;
      RECT 33.339 43.473 35.909 43.529 ;
      RECT 33.385 43.427 35.955 43.483 ;
      RECT 33.431 43.381 36.001 43.437 ;
      RECT 33.477 43.335 36.047 43.391 ;
      RECT 33.523 43.289 36.093 43.345 ;
      RECT 33.569 43.243 36.139 43.299 ;
      RECT 33.615 43.197 36.185 43.253 ;
      RECT 33.661 43.151 36.231 43.207 ;
      RECT 33.707 43.105 36.277 43.161 ;
      RECT 33.753 43.059 36.323 43.115 ;
      RECT 33.799 43.013 36.369 43.069 ;
      RECT 33.845 42.967 36.415 43.023 ;
      RECT 33.891 42.921 36.461 42.977 ;
      RECT 33.937 42.875 36.507 42.931 ;
      RECT 33.983 42.829 36.553 42.885 ;
      RECT 34.029 42.783 36.599 42.839 ;
      RECT 34.075 42.737 36.645 42.793 ;
      RECT 34.121 42.691 36.691 42.747 ;
      RECT 34.167 42.645 36.737 42.701 ;
      RECT 34.213 42.599 36.783 42.655 ;
      RECT 34.259 42.553 36.829 42.609 ;
      RECT 34.305 42.507 36.875 42.563 ;
      RECT 34.351 42.461 36.921 42.517 ;
      RECT 34.397 42.415 36.967 42.471 ;
      RECT 34.443 42.369 37.013 42.425 ;
      RECT 34.489 42.323 37.059 42.379 ;
      RECT 34.535 42.277 37.105 42.333 ;
      RECT 34.581 42.231 37.151 42.287 ;
      RECT 34.627 42.185 37.197 42.241 ;
      RECT 34.673 42.139 37.243 42.195 ;
      RECT 34.719 42.093 37.289 42.149 ;
      RECT 34.765 42.047 37.335 42.103 ;
      RECT 34.811 42.001 37.381 42.057 ;
      RECT 34.857 41.955 37.427 42.011 ;
      RECT 34.903 41.909 37.473 41.965 ;
      RECT 34.949 41.863 37.519 41.919 ;
      RECT 34.995 41.817 37.565 41.873 ;
      RECT 35.041 41.771 37.611 41.827 ;
      RECT 35.087 41.725 37.657 41.781 ;
      RECT 35.133 41.679 37.703 41.735 ;
      RECT 35.179 41.633 37.749 41.689 ;
      RECT 35.225 41.587 37.795 41.643 ;
      RECT 35.271 41.541 37.841 41.597 ;
      RECT 35.317 41.495 37.887 41.551 ;
      RECT 35.363 41.449 37.933 41.505 ;
      RECT 35.409 41.403 37.979 41.459 ;
      RECT 35.455 41.357 38.025 41.413 ;
      RECT 35.501 41.311 38.071 41.367 ;
      RECT 35.547 41.265 38.117 41.321 ;
      RECT 35.593 41.219 38.163 41.275 ;
      RECT 35.639 41.173 38.209 41.229 ;
      RECT 35.685 41.127 38.255 41.183 ;
      RECT 35.731 41.081 38.301 41.137 ;
      RECT 35.777 41.035 38.347 41.091 ;
      RECT 35.823 40.989 38.393 41.045 ;
      RECT 35.869 40.943 38.439 40.999 ;
      RECT 35.915 40.897 38.485 40.953 ;
      RECT 35.961 40.851 38.531 40.907 ;
      RECT 36.007 40.805 38.577 40.861 ;
      RECT 36.053 40.759 38.623 40.815 ;
      RECT 36.099 40.713 38.669 40.769 ;
      RECT 36.145 40.667 38.715 40.723 ;
      RECT 36.191 40.621 38.761 40.677 ;
      RECT 36.237 40.575 38.807 40.631 ;
      RECT 36.283 40.529 38.853 40.585 ;
      RECT 36.329 40.483 38.899 40.539 ;
      RECT 36.375 40.437 38.945 40.493 ;
      RECT 36.421 40.391 38.991 40.447 ;
      RECT 36.467 40.345 39.037 40.401 ;
      RECT 36.513 40.299 39.083 40.355 ;
      RECT 36.559 40.253 39.129 40.309 ;
      RECT 36.605 40.207 39.175 40.263 ;
      RECT 36.651 40.161 39.221 40.217 ;
      RECT 36.697 40.115 39.267 40.171 ;
      RECT 36.743 40.069 39.313 40.125 ;
      RECT 36.789 40.023 39.359 40.079 ;
      RECT 36.835 39.977 39.405 40.033 ;
      RECT 36.881 39.931 39.451 39.987 ;
      RECT 36.927 39.885 39.497 39.941 ;
      RECT 36.973 39.839 39.543 39.895 ;
      RECT 37.019 39.793 39.589 39.849 ;
      RECT 37.065 39.747 39.635 39.803 ;
      RECT 37.111 39.701 39.681 39.757 ;
      RECT 37.157 39.655 39.727 39.711 ;
      RECT 37.203 39.609 39.773 39.665 ;
      RECT 37.249 39.563 39.819 39.619 ;
      RECT 37.295 39.517 39.865 39.573 ;
      RECT 37.341 39.471 39.911 39.527 ;
      RECT 37.387 39.425 39.957 39.481 ;
      RECT 37.433 39.379 40.003 39.435 ;
      RECT 37.479 39.333 40.049 39.389 ;
      RECT 37.525 39.287 40.095 39.343 ;
      RECT 37.571 39.241 40.141 39.297 ;
      RECT 37.617 39.195 40.187 39.251 ;
      RECT 37.663 39.149 40.233 39.205 ;
      RECT 37.709 39.103 40.279 39.159 ;
      RECT 37.755 39.057 40.325 39.113 ;
      RECT 37.801 39.011 40.371 39.067 ;
      RECT 37.847 38.965 40.417 39.021 ;
      RECT 37.893 38.919 40.463 38.975 ;
      RECT 37.939 38.873 40.509 38.929 ;
      RECT 37.985 38.827 40.555 38.883 ;
      RECT 38.031 38.781 40.601 38.837 ;
      RECT 38.077 38.735 40.647 38.791 ;
      RECT 38.123 38.689 40.693 38.745 ;
      RECT 38.169 38.643 40.739 38.699 ;
      RECT 38.215 38.597 40.785 38.653 ;
      RECT 38.261 38.551 40.831 38.607 ;
      RECT 38.307 38.505 40.877 38.561 ;
      RECT 38.353 38.459 40.923 38.515 ;
      RECT 38.399 38.413 40.969 38.469 ;
      RECT 38.445 38.367 41.015 38.423 ;
      RECT 38.491 38.321 41.061 38.377 ;
      RECT 38.537 38.275 41.107 38.331 ;
      RECT 38.583 38.229 41.153 38.285 ;
      RECT 38.629 38.183 41.199 38.239 ;
      RECT 38.675 38.137 41.245 38.193 ;
      RECT 38.721 38.091 41.291 38.147 ;
      RECT 38.767 38.045 41.337 38.101 ;
      RECT 38.813 37.999 41.383 38.055 ;
      RECT 38.859 37.953 41.429 38.009 ;
      RECT 38.905 37.907 41.475 37.963 ;
      RECT 38.951 37.861 41.521 37.917 ;
      RECT 38.997 37.815 41.567 37.871 ;
      RECT 39.043 37.769 41.613 37.825 ;
      RECT 39.089 37.723 41.659 37.779 ;
      RECT 39.135 37.677 41.705 37.733 ;
      RECT 39.181 37.631 41.751 37.687 ;
      RECT 39.227 37.585 41.797 37.641 ;
      RECT 39.273 37.539 41.843 37.595 ;
      RECT 39.319 37.493 41.889 37.549 ;
      RECT 39.365 37.447 41.935 37.503 ;
      RECT 39.411 37.401 41.981 37.457 ;
      RECT 39.457 37.355 42.027 37.411 ;
      RECT 39.503 37.309 42.073 37.365 ;
      RECT 39.549 37.263 42.119 37.319 ;
      RECT 39.595 37.217 42.165 37.273 ;
      RECT 39.641 37.171 42.211 37.227 ;
      RECT 39.687 37.125 42.257 37.181 ;
      RECT 39.733 37.079 42.303 37.135 ;
      RECT 39.779 37.033 42.349 37.089 ;
      RECT 39.825 36.987 42.395 37.043 ;
      RECT 39.871 36.941 42.441 36.997 ;
      RECT 39.917 36.895 42.487 36.951 ;
      RECT 39.963 36.849 42.533 36.905 ;
      RECT 40.009 36.803 42.579 36.859 ;
      RECT 40.055 36.757 42.625 36.813 ;
      RECT 40.101 36.711 42.671 36.767 ;
      RECT 40.147 36.665 42.717 36.721 ;
      RECT 40.193 36.619 42.763 36.675 ;
      RECT 40.239 36.573 42.809 36.629 ;
      RECT 40.285 36.527 42.855 36.583 ;
      RECT 40.331 36.481 42.901 36.537 ;
      RECT 40.377 36.435 42.947 36.491 ;
      RECT 40.423 36.389 42.993 36.445 ;
      RECT 40.469 36.343 43.039 36.399 ;
      RECT 40.515 36.297 43.085 36.353 ;
      RECT 40.561 36.251 43.131 36.307 ;
      RECT 40.607 36.205 43.177 36.261 ;
      RECT 40.653 36.159 43.223 36.215 ;
      RECT 40.699 36.113 43.269 36.169 ;
      RECT 40.745 36.067 43.315 36.123 ;
      RECT 40.791 36.021 43.361 36.077 ;
      RECT 40.837 35.975 43.407 36.031 ;
      RECT 40.883 35.929 43.453 35.985 ;
      RECT 40.929 35.883 43.499 35.939 ;
      RECT 40.975 35.837 43.545 35.893 ;
      RECT 41.021 35.791 43.591 35.847 ;
      RECT 41.067 35.745 43.637 35.801 ;
      RECT 41.113 35.699 43.683 35.755 ;
      RECT 41.159 35.653 43.729 35.709 ;
      RECT 41.205 35.607 43.775 35.663 ;
      RECT 41.251 35.561 43.821 35.617 ;
      RECT 41.297 35.515 43.867 35.571 ;
      RECT 41.343 35.469 43.913 35.525 ;
      RECT 41.389 35.423 43.959 35.479 ;
      RECT 41.435 35.377 44.005 35.433 ;
      RECT 41.481 35.331 44.051 35.387 ;
      RECT 41.527 35.285 44.097 35.341 ;
      RECT 41.573 35.239 44.143 35.295 ;
      RECT 41.619 35.193 44.189 35.249 ;
      RECT 41.665 35.147 44.235 35.203 ;
      RECT 41.711 35.101 44.281 35.157 ;
      RECT 41.757 35.055 44.327 35.111 ;
      RECT 41.803 35.009 44.373 35.065 ;
      RECT 41.849 34.963 44.419 35.019 ;
      RECT 41.895 34.917 44.465 34.973 ;
      RECT 41.941 34.871 44.511 34.927 ;
      RECT 41.987 34.825 44.557 34.881 ;
      RECT 42.033 34.779 44.603 34.835 ;
      RECT 42.079 34.733 44.649 34.789 ;
      RECT 42.125 34.687 44.695 34.743 ;
      RECT 42.171 34.641 44.741 34.697 ;
      RECT 42.217 34.595 44.787 34.651 ;
      RECT 42.263 34.549 44.833 34.605 ;
      RECT 42.309 34.503 44.879 34.559 ;
      RECT 42.355 34.457 44.925 34.513 ;
      RECT 42.401 34.411 44.971 34.467 ;
      RECT 42.447 34.365 45.017 34.421 ;
      RECT 42.493 34.319 45.063 34.375 ;
      RECT 42.539 34.273 45.109 34.329 ;
      RECT 42.585 34.227 45.155 34.283 ;
      RECT 42.631 34.181 45.201 34.237 ;
      RECT 42.677 34.135 45.247 34.191 ;
      RECT 42.723 34.089 45.293 34.145 ;
      RECT 42.769 34.043 45.339 34.099 ;
      RECT 42.815 33.997 45.385 34.053 ;
      RECT 42.861 33.951 45.431 34.007 ;
      RECT 42.907 33.905 45.477 33.961 ;
      RECT 42.953 33.859 45.523 33.915 ;
      RECT 42.999 33.813 45.569 33.869 ;
      RECT 43.045 33.767 45.615 33.823 ;
      RECT 43.091 33.721 45.661 33.777 ;
      RECT 43.137 33.675 45.707 33.731 ;
      RECT 43.183 33.629 45.753 33.685 ;
      RECT 43.229 33.583 45.799 33.639 ;
      RECT 43.275 33.537 45.845 33.593 ;
      RECT 43.321 33.491 45.891 33.547 ;
      RECT 43.367 33.445 45.937 33.501 ;
      RECT 43.413 33.399 45.983 33.455 ;
      RECT 43.459 33.353 46.029 33.409 ;
      RECT 43.505 33.307 46.075 33.363 ;
      RECT 43.551 33.261 46.121 33.317 ;
      RECT 43.597 33.215 46.167 33.271 ;
      RECT 43.643 33.169 46.213 33.225 ;
      RECT 43.689 33.123 46.259 33.179 ;
      RECT 43.735 33.077 46.305 33.133 ;
      RECT 43.781 33.031 46.351 33.087 ;
      RECT 43.827 32.985 46.397 33.041 ;
      RECT 43.873 32.939 46.443 32.995 ;
      RECT 43.919 32.893 46.489 32.949 ;
      RECT 43.965 32.847 46.535 32.903 ;
      RECT 44.011 32.801 46.581 32.857 ;
      RECT 44.057 32.755 46.627 32.811 ;
      RECT 44.103 32.709 46.673 32.765 ;
      RECT 44.149 32.663 46.719 32.719 ;
      RECT 44.195 32.617 46.765 32.673 ;
      RECT 44.241 32.571 46.811 32.627 ;
      RECT 44.287 32.525 46.857 32.581 ;
      RECT 44.333 32.479 46.903 32.535 ;
      RECT 44.379 32.433 46.949 32.489 ;
      RECT 44.425 32.387 46.995 32.443 ;
      RECT 44.471 32.341 47.041 32.397 ;
      RECT 44.517 32.295 47.087 32.351 ;
      RECT 44.563 32.249 47.133 32.305 ;
      RECT 44.609 32.203 47.179 32.259 ;
      RECT 44.655 32.157 47.225 32.213 ;
      RECT 44.701 32.111 47.271 32.167 ;
      RECT 44.747 32.065 47.317 32.121 ;
      RECT 44.793 32.019 47.363 32.075 ;
      RECT 44.839 31.973 47.409 32.029 ;
      RECT 44.885 31.927 47.455 31.983 ;
      RECT 44.931 31.881 47.501 31.937 ;
      RECT 44.977 31.835 47.547 31.891 ;
      RECT 45.023 31.789 47.593 31.845 ;
      RECT 45.069 31.743 47.639 31.799 ;
      RECT 45.115 31.697 47.685 31.753 ;
      RECT 45.161 31.651 47.731 31.707 ;
      RECT 45.207 31.605 47.777 31.661 ;
      RECT 45.253 31.559 47.823 31.615 ;
      RECT 45.299 31.513 47.869 31.569 ;
      RECT 45.345 31.467 47.915 31.523 ;
      RECT 45.391 31.421 47.961 31.477 ;
      RECT 45.437 31.375 48.007 31.431 ;
      RECT 45.483 31.329 48.053 31.385 ;
      RECT 45.529 31.283 48.099 31.339 ;
      RECT 45.575 31.237 48.145 31.293 ;
      RECT 45.621 31.191 48.191 31.247 ;
      RECT 45.667 31.145 48.237 31.201 ;
      RECT 45.713 31.099 48.283 31.155 ;
      RECT 45.759 31.053 48.329 31.109 ;
      RECT 45.805 31.007 48.375 31.063 ;
      RECT 45.851 30.961 48.421 31.017 ;
      RECT 45.897 30.915 48.467 30.971 ;
      RECT 45.943 30.869 48.513 30.925 ;
      RECT 45.989 30.823 48.559 30.879 ;
      RECT 46.035 30.777 48.605 30.833 ;
      RECT 46.081 30.731 48.651 30.787 ;
      RECT 46.127 30.685 48.697 30.741 ;
      RECT 46.173 30.639 48.743 30.695 ;
      RECT 46.219 30.593 48.789 30.649 ;
      RECT 46.265 30.547 48.835 30.603 ;
      RECT 46.311 30.501 48.881 30.557 ;
      RECT 46.357 30.455 48.927 30.511 ;
      RECT 46.403 30.409 48.973 30.465 ;
      RECT 46.449 30.363 49.019 30.419 ;
      RECT 46.495 30.317 49.065 30.373 ;
      RECT 46.541 30.271 49.111 30.327 ;
      RECT 46.587 30.225 49.157 30.281 ;
      RECT 46.633 30.179 49.203 30.235 ;
      RECT 46.679 30.133 49.249 30.189 ;
      RECT 46.725 30.087 49.295 30.143 ;
      RECT 46.771 30.041 49.341 30.097 ;
      RECT 46.817 29.995 49.387 30.051 ;
      RECT 46.863 29.949 49.433 30.005 ;
      RECT 46.909 29.903 49.479 29.959 ;
      RECT 46.955 29.857 49.525 29.913 ;
      RECT 47.001 29.811 49.571 29.867 ;
      RECT 47.047 29.765 49.617 29.821 ;
      RECT 47.093 29.719 49.663 29.775 ;
      RECT 47.139 29.673 49.709 29.729 ;
      RECT 47.185 29.627 49.755 29.683 ;
      RECT 47.231 29.581 49.801 29.637 ;
      RECT 47.277 29.535 49.847 29.591 ;
      RECT 47.323 29.489 49.893 29.545 ;
      RECT 47.369 29.443 49.939 29.499 ;
      RECT 47.415 29.397 49.985 29.453 ;
      RECT 47.461 29.351 50.031 29.407 ;
      RECT 47.507 29.305 50.077 29.361 ;
      RECT 47.553 29.259 50.123 29.315 ;
      RECT 47.599 29.213 50.169 29.269 ;
      RECT 47.645 29.167 50.215 29.223 ;
      RECT 47.691 29.121 50.261 29.177 ;
      RECT 47.737 29.075 50.307 29.131 ;
      RECT 47.783 29.029 50.353 29.085 ;
      RECT 47.829 28.983 50.399 29.039 ;
      RECT 47.875 28.937 50.445 28.993 ;
      RECT 47.921 28.891 50.491 28.947 ;
      RECT 47.967 28.845 50.537 28.901 ;
      RECT 48.013 28.799 50.583 28.855 ;
      RECT 48.059 28.753 50.629 28.809 ;
      RECT 48.105 28.707 50.675 28.763 ;
      RECT 48.151 28.661 50.721 28.717 ;
      RECT 48.197 28.615 50.767 28.671 ;
      RECT 48.243 28.569 50.813 28.625 ;
      RECT 48.289 28.523 50.859 28.579 ;
      RECT 48.335 28.477 50.905 28.533 ;
      RECT 48.381 28.431 50.951 28.487 ;
      RECT 48.427 28.385 50.997 28.441 ;
      RECT 48.473 28.339 51.043 28.395 ;
      RECT 48.519 28.293 51.089 28.349 ;
      RECT 48.565 28.247 51.135 28.303 ;
      RECT 48.611 28.201 51.181 28.257 ;
      RECT 48.657 28.155 51.227 28.211 ;
      RECT 48.703 28.109 51.273 28.165 ;
      RECT 48.749 28.063 51.319 28.119 ;
      RECT 48.795 28.017 51.365 28.073 ;
      RECT 48.841 27.971 51.411 28.027 ;
      RECT 48.887 27.925 51.457 27.981 ;
      RECT 48.933 27.879 51.503 27.935 ;
      RECT 48.979 27.833 51.549 27.889 ;
      RECT 49.025 27.787 51.595 27.843 ;
      RECT 49.071 27.741 51.641 27.797 ;
      RECT 49.117 27.695 51.687 27.751 ;
      RECT 49.163 27.649 51.733 27.705 ;
      RECT 49.209 27.603 51.779 27.659 ;
      RECT 49.255 27.557 51.825 27.613 ;
      RECT 49.301 27.511 51.871 27.567 ;
      RECT 49.347 27.465 51.917 27.521 ;
      RECT 49.393 27.419 51.963 27.475 ;
      RECT 49.439 27.373 52.009 27.429 ;
      RECT 49.485 27.327 52.055 27.383 ;
      RECT 49.531 27.281 52.101 27.337 ;
      RECT 49.577 27.235 52.147 27.291 ;
      RECT 49.623 27.189 52.193 27.245 ;
      RECT 49.669 27.143 52.239 27.199 ;
      RECT 49.715 27.097 52.285 27.153 ;
      RECT 49.761 27.051 52.331 27.107 ;
      RECT 49.807 27.005 52.377 27.061 ;
      RECT 49.853 26.959 52.423 27.015 ;
      RECT 49.899 26.913 52.469 26.969 ;
      RECT 49.945 26.867 52.515 26.923 ;
      RECT 49.991 26.821 52.561 26.877 ;
      RECT 50.037 26.775 52.607 26.831 ;
      RECT 50.083 26.729 52.653 26.785 ;
      RECT 50.129 26.683 52.699 26.739 ;
      RECT 50.175 26.637 52.745 26.693 ;
      RECT 50.221 26.591 52.791 26.647 ;
      RECT 50.267 26.545 52.837 26.601 ;
      RECT 50.313 26.499 52.883 26.555 ;
      RECT 50.359 26.453 52.929 26.509 ;
      RECT 50.405 26.407 52.975 26.463 ;
      RECT 50.451 26.361 53.021 26.417 ;
      RECT 50.497 26.315 53.067 26.371 ;
      RECT 50.543 26.269 53.113 26.325 ;
      RECT 50.589 26.223 53.159 26.279 ;
      RECT 50.635 26.177 53.205 26.233 ;
      RECT 50.681 26.131 53.251 26.187 ;
      RECT 50.727 26.085 53.297 26.141 ;
      RECT 50.773 26.039 53.343 26.095 ;
      RECT 50.819 25.993 53.389 26.049 ;
      RECT 50.865 25.947 53.435 26.003 ;
      RECT 50.911 25.901 53.481 25.957 ;
      RECT 50.957 25.855 53.527 25.911 ;
      RECT 51.003 25.809 53.573 25.865 ;
      RECT 51.049 25.763 53.619 25.819 ;
      RECT 51.095 25.717 53.665 25.773 ;
      RECT 51.141 25.671 53.711 25.727 ;
      RECT 51.187 25.625 53.757 25.681 ;
      RECT 51.233 25.579 53.803 25.635 ;
      RECT 51.279 25.533 53.849 25.589 ;
      RECT 51.325 25.487 53.895 25.543 ;
      RECT 51.371 25.441 53.941 25.497 ;
      RECT 51.417 25.395 53.987 25.451 ;
      RECT 51.463 25.349 54.033 25.405 ;
      RECT 51.509 25.303 54.079 25.359 ;
      RECT 51.555 25.257 54.125 25.313 ;
      RECT 51.601 25.211 54.171 25.267 ;
      RECT 51.647 25.165 54.217 25.221 ;
      RECT 51.693 25.119 54.263 25.175 ;
      RECT 51.739 25.073 54.309 25.129 ;
      RECT 51.785 25.027 54.355 25.083 ;
      RECT 51.831 24.981 54.401 25.037 ;
      RECT 51.877 24.935 54.447 24.991 ;
      RECT 51.923 24.889 54.493 24.945 ;
      RECT 51.969 24.843 54.539 24.899 ;
      RECT 52.015 24.797 54.585 24.853 ;
      RECT 52.061 24.751 54.631 24.807 ;
      RECT 52.107 24.705 54.677 24.761 ;
      RECT 52.153 24.659 54.723 24.715 ;
      RECT 52.199 24.613 54.769 24.669 ;
      RECT 52.245 24.567 54.815 24.623 ;
      RECT 52.291 24.521 54.861 24.577 ;
      RECT 52.337 24.475 54.907 24.531 ;
      RECT 52.383 24.429 54.953 24.485 ;
      RECT 52.429 24.383 54.999 24.439 ;
      RECT 52.475 24.337 55.045 24.393 ;
      RECT 52.521 24.291 55.091 24.347 ;
      RECT 52.567 24.245 55.137 24.301 ;
      RECT 52.613 24.199 55.183 24.255 ;
      RECT 52.659 24.153 55.229 24.209 ;
      RECT 52.705 24.107 55.275 24.163 ;
      RECT 52.751 24.061 55.321 24.117 ;
      RECT 52.797 24.015 55.367 24.071 ;
      RECT 52.843 23.969 55.413 24.025 ;
      RECT 52.889 23.923 55.459 23.979 ;
      RECT 52.935 23.877 55.505 23.933 ;
      RECT 52.981 23.831 55.551 23.887 ;
      RECT 53.027 23.785 55.597 23.841 ;
      RECT 53.073 23.739 55.643 23.795 ;
      RECT 53.119 23.693 55.689 23.749 ;
      RECT 53.165 23.647 55.735 23.703 ;
      RECT 53.211 23.601 55.781 23.657 ;
      RECT 53.257 23.555 55.827 23.611 ;
      RECT 53.303 23.509 55.873 23.565 ;
      RECT 53.349 23.463 55.919 23.519 ;
      RECT 53.395 23.417 55.965 23.473 ;
      RECT 53.441 23.371 56.011 23.427 ;
      RECT 53.487 23.325 56.057 23.381 ;
      RECT 53.533 23.279 56.103 23.335 ;
      RECT 53.579 23.233 56.149 23.289 ;
      RECT 53.625 23.187 56.195 23.243 ;
      RECT 53.671 23.141 56.241 23.197 ;
      RECT 53.717 23.095 56.287 23.151 ;
      RECT 53.763 23.049 56.333 23.105 ;
      RECT 53.809 23.003 56.379 23.059 ;
      RECT 53.855 22.957 56.425 23.013 ;
      RECT 53.901 22.911 56.471 22.967 ;
      RECT 53.947 22.865 56.517 22.921 ;
      RECT 53.993 22.819 56.563 22.875 ;
      RECT 54.039 22.773 56.609 22.829 ;
      RECT 54.085 22.727 56.655 22.783 ;
      RECT 54.131 22.681 56.701 22.737 ;
      RECT 54.177 22.635 56.747 22.691 ;
      RECT 54.223 22.589 56.793 22.645 ;
      RECT 54.269 22.543 56.839 22.599 ;
      RECT 54.315 22.497 56.885 22.553 ;
      RECT 54.361 22.451 56.931 22.507 ;
      RECT 54.407 22.405 56.977 22.461 ;
      RECT 54.453 22.359 57.023 22.415 ;
      RECT 54.499 22.313 57.069 22.369 ;
      RECT 54.545 22.267 57.115 22.323 ;
      RECT 54.591 22.221 57.161 22.277 ;
      RECT 54.637 22.175 57.207 22.231 ;
      RECT 54.683 22.129 57.253 22.185 ;
      RECT 54.729 22.083 57.299 22.139 ;
      RECT 54.775 22.037 57.345 22.093 ;
      RECT 54.821 21.991 57.391 22.047 ;
      RECT 54.867 21.945 57.437 22.001 ;
      RECT 54.913 21.899 57.483 21.955 ;
      RECT 54.959 21.853 57.529 21.909 ;
      RECT 55.005 21.807 57.575 21.863 ;
      RECT 55.051 21.761 57.621 21.817 ;
      RECT 55.097 21.715 57.667 21.771 ;
      RECT 55.143 21.669 57.713 21.725 ;
      RECT 55.189 21.623 57.759 21.679 ;
      RECT 55.235 21.577 57.805 21.633 ;
      RECT 55.281 21.531 57.851 21.587 ;
      RECT 55.327 21.485 57.897 21.541 ;
      RECT 55.373 21.439 57.943 21.495 ;
      RECT 55.419 21.393 57.989 21.449 ;
      RECT 55.465 21.347 58.035 21.403 ;
      RECT 55.511 21.301 58.081 21.357 ;
      RECT 55.557 21.255 58.127 21.311 ;
      RECT 55.603 21.209 58.173 21.265 ;
      RECT 55.649 21.163 58.219 21.219 ;
      RECT 55.695 21.117 58.265 21.173 ;
      RECT 55.741 21.071 58.311 21.127 ;
      RECT 55.787 21.025 58.357 21.081 ;
      RECT 55.833 20.979 58.403 21.035 ;
      RECT 55.879 20.933 58.449 20.989 ;
      RECT 55.925 20.887 58.495 20.943 ;
      RECT 55.971 20.841 58.541 20.897 ;
      RECT 56.017 20.795 58.587 20.851 ;
      RECT 56.063 20.749 58.633 20.805 ;
      RECT 56.109 20.703 58.679 20.759 ;
      RECT 56.155 20.663 58.725 20.713 ;
      RECT 56.19 20.622 58.771 20.667 ;
      RECT 56.236 20.576 58.817 20.621 ;
      RECT 56.282 20.53 58.863 20.575 ;
      RECT 56.328 20.484 58.909 20.529 ;
      RECT 56.374 20.438 58.955 20.483 ;
      RECT 56.42 20.392 59.001 20.437 ;
      RECT 56.466 20.346 59.047 20.391 ;
      RECT 56.512 20.3 59.093 20.345 ;
      RECT 56.558 20.254 59.139 20.299 ;
      RECT 56.604 20.208 59.185 20.253 ;
      RECT 56.65 20.162 59.231 20.207 ;
      RECT 56.696 20.116 59.277 20.161 ;
      RECT 56.742 20.07 59.323 20.115 ;
      RECT 56.788 20.024 59.369 20.069 ;
      RECT 56.834 19.978 59.415 20.023 ;
      RECT 56.88 19.932 59.461 19.977 ;
      RECT 56.926 19.886 59.507 19.931 ;
      RECT 56.972 19.84 59.553 19.885 ;
      RECT 57.018 19.794 59.599 19.839 ;
      RECT 57.064 19.748 59.645 19.793 ;
      RECT 57.11 19.702 59.691 19.747 ;
      RECT 57.156 19.656 59.737 19.701 ;
      RECT 57.202 19.61 59.783 19.655 ;
      RECT 57.248 19.564 59.829 19.609 ;
      RECT 57.294 19.518 59.875 19.563 ;
      RECT 57.34 19.472 59.921 19.517 ;
      RECT 57.386 19.426 59.967 19.471 ;
      RECT 57.432 19.38 60.013 19.425 ;
      RECT 57.478 19.334 60.059 19.379 ;
      RECT 57.524 19.288 60.105 19.333 ;
      RECT 57.57 19.242 60.151 19.287 ;
      RECT 57.616 19.196 60.197 19.241 ;
      RECT 57.662 19.15 60.243 19.195 ;
      RECT 57.708 19.104 60.289 19.149 ;
      RECT 57.754 19.058 60.335 19.103 ;
      RECT 57.8 19.012 60.381 19.057 ;
      RECT 57.846 18.966 60.427 19.011 ;
      RECT 57.892 18.92 60.473 18.965 ;
      RECT 57.938 18.874 60.519 18.919 ;
      RECT 57.984 18.828 60.565 18.873 ;
      RECT 58.03 18.782 60.611 18.827 ;
      RECT 58.076 18.736 60.657 18.781 ;
      RECT 58.122 18.69 60.703 18.735 ;
      RECT 58.168 18.644 60.749 18.689 ;
      RECT 58.214 18.598 60.795 18.643 ;
      RECT 58.26 18.552 60.841 18.597 ;
      RECT 58.306 18.506 60.887 18.551 ;
      RECT 58.352 18.46 60.933 18.505 ;
      RECT 58.398 18.414 60.979 18.459 ;
      RECT 58.444 18.368 61.025 18.413 ;
      RECT 58.49 18.322 61.071 18.367 ;
      RECT 58.536 18.276 61.117 18.321 ;
      RECT 58.582 18.23 61.163 18.275 ;
      RECT 58.628 18.184 61.209 18.229 ;
      RECT 58.674 18.138 61.255 18.183 ;
      RECT 58.72 18.092 61.301 18.137 ;
      RECT 58.766 18.046 61.347 18.091 ;
      RECT 58.812 18 61.393 18.045 ;
      RECT 58.858 17.954 61.439 17.999 ;
      RECT 58.904 17.908 61.485 17.953 ;
      RECT 58.95 17.862 61.531 17.907 ;
      RECT 58.996 17.816 61.577 17.861 ;
      RECT 59.042 17.77 61.623 17.815 ;
      RECT 59.088 17.724 61.669 17.769 ;
      RECT 59.134 17.678 61.715 17.723 ;
      RECT 59.18 17.632 61.761 17.677 ;
      RECT 59.226 17.586 61.807 17.631 ;
      RECT 59.272 17.54 61.853 17.585 ;
      RECT 59.318 17.494 61.899 17.539 ;
      RECT 59.364 17.448 61.945 17.493 ;
      RECT 59.41 17.402 61.991 17.447 ;
      RECT 59.456 17.356 62.037 17.401 ;
      RECT 59.502 17.31 62.083 17.355 ;
      RECT 59.548 17.264 62.129 17.309 ;
      RECT 59.594 17.218 62.175 17.263 ;
      RECT 59.64 17.172 62.221 17.217 ;
      RECT 59.686 17.126 62.267 17.171 ;
      RECT 59.732 17.08 62.313 17.125 ;
      RECT 59.778 17.034 62.359 17.079 ;
      RECT 59.824 16.988 62.405 17.033 ;
      RECT 59.87 16.942 62.451 16.987 ;
      RECT 59.916 16.896 62.497 16.941 ;
      RECT 59.962 16.85 62.543 16.895 ;
      RECT 60.008 16.804 62.589 16.849 ;
      RECT 61.158 15.675 110 16.825 ;
      RECT 60.054 16.758 110 16.825 ;
      RECT 61.112 15.699 61.163 18.275 ;
      RECT 60.1 16.712 110 16.825 ;
      RECT 61.066 15.746 61.117 18.321 ;
      RECT 60.146 16.666 110 16.825 ;
      RECT 61.02 15.792 61.071 18.367 ;
      RECT 60.192 16.62 110 16.825 ;
      RECT 60.974 15.838 61.025 18.413 ;
      RECT 60.238 16.574 110 16.825 ;
      RECT 60.928 15.884 60.979 18.459 ;
      RECT 60.284 16.528 110 16.825 ;
      RECT 60.882 15.93 60.933 18.505 ;
      RECT 60.33 16.482 110 16.825 ;
      RECT 60.836 15.976 60.887 18.551 ;
      RECT 60.376 16.436 110 16.825 ;
      RECT 60.79 16.022 60.841 18.597 ;
      RECT 60.422 16.39 110 16.825 ;
      RECT 60.744 16.068 60.795 18.643 ;
      RECT 60.468 16.344 110 16.825 ;
      RECT 60.698 16.114 60.749 18.689 ;
      RECT 60.514 16.298 110 16.825 ;
      RECT 60.652 16.16 60.703 18.735 ;
      RECT 60.56 16.252 110 16.825 ;
      RECT 60.606 16.206 60.657 18.781 ;
      RECT 29.175 67.887 30.325 110 ;
      RECT 29.175 67.887 30.371 69.317 ;
      RECT 29.175 67.887 30.417 69.271 ;
      RECT 29.175 67.887 30.463 69.225 ;
      RECT 29.175 67.887 30.509 69.179 ;
      RECT 29.175 67.887 30.555 69.133 ;
      RECT 29.175 67.887 30.601 69.087 ;
      RECT 29.175 67.887 30.647 69.041 ;
      RECT 29.175 67.887 30.693 68.995 ;
      RECT 29.175 67.887 30.739 68.949 ;
      RECT 29.175 67.887 30.785 68.903 ;
      RECT 29.175 67.887 30.831 68.857 ;
      RECT 29.175 67.887 30.877 68.811 ;
      RECT 29.175 67.887 30.923 68.765 ;
      RECT 29.175 67.887 30.969 68.719 ;
      RECT 29.175 67.887 31.015 68.673 ;
      RECT 29.175 67.887 31.061 68.627 ;
      RECT 29.175 67.887 31.107 68.581 ;
      RECT 29.175 67.887 31.153 68.535 ;
      RECT 29.175 67.887 31.199 68.489 ;
      RECT 29.175 67.887 31.245 68.443 ;
      RECT 29.175 67.887 31.291 68.397 ;
      RECT 29.175 67.887 31.337 68.351 ;
      RECT 29.175 67.887 31.383 68.305 ;
      RECT 29.175 67.887 31.429 68.259 ;
      RECT 29.175 67.887 31.475 68.213 ;
      RECT 29.175 67.887 31.521 68.167 ;
      RECT 29.175 67.887 31.567 68.121 ;
      RECT 29.175 67.887 31.613 68.075 ;
      RECT 29.175 67.887 31.659 68.029 ;
      RECT 29.175 67.887 31.705 67.983 ;
      RECT 29.175 67.887 31.751 67.937 ;
      RECT 29.221 67.841 31.797 67.891 ;
      RECT 29.267 67.795 31.843 67.845 ;
      RECT 29.313 67.749 31.889 67.799 ;
      RECT 29.359 67.703 31.935 67.753 ;
      RECT 29.405 67.657 31.981 67.707 ;
      RECT 29.451 67.611 32.027 67.661 ;
      RECT 29.497 67.565 32.073 67.615 ;
      RECT 29.543 67.519 32.119 67.569 ;
      RECT 29.589 67.473 32.165 67.523 ;
      RECT 29.635 67.427 32.211 67.477 ;
      RECT 29.681 67.381 32.257 67.431 ;
      RECT 29.727 67.335 32.303 67.385 ;
      RECT 29.773 67.289 32.349 67.339 ;
      RECT 29.819 67.243 32.395 67.293 ;
      RECT 29.865 67.197 32.441 67.247 ;
      RECT 29.911 67.151 32.487 67.201 ;
      RECT 29.957 67.105 32.533 67.155 ;
      RECT 30.003 67.059 32.579 67.109 ;
      RECT 30.049 67.013 32.625 67.063 ;
      RECT 30.095 66.967 32.671 67.017 ;
      RECT 30.141 66.921 32.717 66.971 ;
      RECT 30.187 66.875 32.763 66.925 ;
      RECT 30.233 66.829 32.809 66.879 ;
      RECT 30.279 66.783 32.855 66.833 ;
      RECT 30.325 66.737 32.901 66.787 ;
      RECT 30.371 66.691 32.947 66.741 ;
      RECT 30.417 66.645 32.993 66.695 ;
      RECT 30.463 66.599 33.039 66.649 ;
      RECT 30.509 66.553 33.085 66.603 ;
      RECT 30.555 66.507 33.131 66.557 ;
      RECT 30.601 66.461 33.177 66.511 ;
      RECT 30.647 66.415 33.223 66.465 ;
      RECT 30.693 66.369 33.269 66.419 ;
      RECT 30.739 66.323 33.315 66.373 ;
      RECT 30.785 66.277 33.361 66.327 ;
      RECT 30.831 66.231 33.407 66.281 ;
      RECT 30.877 66.185 33.453 66.235 ;
      RECT 30.923 66.139 33.499 66.189 ;
      RECT 30.969 66.093 33.545 66.143 ;
      RECT 31.015 66.047 33.591 66.097 ;
      RECT 31.061 66.001 33.637 66.051 ;
      RECT 31.107 65.955 33.683 66.005 ;
      RECT 31.153 65.909 33.729 65.959 ;
      RECT 31.199 65.863 33.775 65.913 ;
      RECT 31.245 65.817 33.821 65.867 ;
      RECT 31.291 65.771 33.867 65.821 ;
      RECT 31.337 65.725 33.913 65.775 ;
      RECT 31.383 65.679 33.959 65.729 ;
      RECT 31.429 65.633 34.005 65.683 ;
      RECT 31.475 65.587 34.051 65.637 ;
      RECT 31.521 65.541 34.097 65.591 ;
      RECT 31.567 65.495 34.143 65.545 ;
      RECT 31.613 65.449 34.189 65.499 ;
      RECT 31.659 65.403 34.235 65.453 ;
      RECT 31.705 65.357 34.281 65.407 ;
      RECT 31.751 65.311 34.327 65.361 ;
      RECT 31.797 65.265 34.373 65.315 ;
      RECT 31.843 65.219 34.419 65.269 ;
      RECT 31.889 65.173 34.465 65.223 ;
      RECT 31.935 65.127 34.511 65.177 ;
      RECT 31.981 65.081 34.557 65.131 ;
      RECT 32.027 65.035 34.603 65.085 ;
      RECT 32.073 64.989 34.649 65.039 ;
      RECT 32.119 64.943 34.695 64.993 ;
      RECT 32.165 64.897 34.741 64.947 ;
      RECT 32.211 64.851 34.787 64.901 ;
      RECT 32.257 64.805 34.833 64.855 ;
      RECT 32.303 64.759 34.879 64.809 ;
      RECT 32.349 64.713 34.925 64.763 ;
      RECT 32.395 64.667 34.971 64.717 ;
      RECT 32.441 64.621 35.017 64.671 ;
      RECT 32.487 64.575 35.063 64.625 ;
      RECT 32.533 64.529 35.109 64.579 ;
      RECT 32.579 64.483 35.155 64.533 ;
      RECT 32.625 64.437 35.201 64.487 ;
      RECT 32.671 64.391 35.247 64.441 ;
      RECT 32.717 64.345 35.293 64.395 ;
      RECT 32.763 64.299 35.339 64.349 ;
      RECT 32.809 64.253 35.385 64.303 ;
      RECT 32.855 64.207 35.431 64.257 ;
      RECT 32.901 64.161 35.477 64.211 ;
      RECT 32.947 64.115 35.523 64.165 ;
      RECT 32.993 64.069 35.569 64.119 ;
      RECT 33.039 64.023 35.615 64.073 ;
      RECT 33.085 63.977 35.661 64.027 ;
      RECT 33.131 63.931 35.707 63.981 ;
      RECT 33.177 63.885 35.753 63.935 ;
      RECT 33.223 63.839 35.799 63.889 ;
      RECT 33.269 63.793 35.845 63.843 ;
      RECT 33.315 63.747 35.891 63.797 ;
      RECT 33.361 63.701 35.937 63.751 ;
      RECT 33.407 63.655 35.983 63.705 ;
      RECT 33.453 63.609 36.029 63.659 ;
      RECT 33.499 63.563 36.075 63.613 ;
      RECT 33.545 63.517 36.121 63.567 ;
      RECT 33.591 63.471 36.167 63.521 ;
      RECT 33.637 63.425 36.213 63.475 ;
      RECT 33.683 63.379 36.259 63.429 ;
      RECT 33.729 63.333 36.305 63.383 ;
      RECT 33.775 63.287 36.351 63.337 ;
      RECT 33.821 63.241 36.397 63.291 ;
      RECT 33.867 63.195 36.443 63.245 ;
      RECT 33.913 63.149 36.489 63.199 ;
      RECT 33.959 63.103 36.535 63.153 ;
      RECT 34.005 63.057 36.581 63.107 ;
      RECT 34.051 63.011 36.627 63.061 ;
      RECT 34.097 62.965 36.673 63.015 ;
      RECT 34.143 62.919 36.719 62.969 ;
      RECT 34.189 62.873 36.765 62.923 ;
      RECT 34.235 62.827 36.811 62.877 ;
      RECT 34.281 62.781 36.857 62.831 ;
      RECT 34.327 62.735 36.903 62.785 ;
      RECT 34.373 62.689 36.949 62.739 ;
      RECT 34.419 62.643 36.995 62.693 ;
      RECT 34.465 62.597 37.041 62.647 ;
      RECT 34.511 62.551 37.087 62.601 ;
      RECT 34.557 62.505 37.133 62.555 ;
      RECT 34.603 62.459 37.179 62.509 ;
      RECT 34.649 62.413 37.225 62.463 ;
      RECT 34.695 62.367 37.271 62.417 ;
      RECT 34.741 62.321 37.317 62.371 ;
      RECT 34.787 62.275 37.363 62.325 ;
      RECT 34.833 62.229 37.409 62.279 ;
      RECT 34.879 62.183 37.455 62.233 ;
      RECT 34.925 62.137 37.501 62.187 ;
      RECT 34.971 62.091 37.547 62.141 ;
      RECT 35.017 62.045 37.593 62.095 ;
      RECT 35.063 61.999 37.639 62.049 ;
      RECT 35.109 61.953 37.685 62.003 ;
      RECT 35.155 61.907 37.731 61.957 ;
      RECT 35.201 61.861 37.777 61.911 ;
      RECT 35.247 61.815 37.823 61.865 ;
      RECT 35.293 61.769 37.869 61.819 ;
      RECT 35.339 61.723 37.915 61.773 ;
      RECT 35.385 61.677 37.961 61.727 ;
      RECT 35.431 61.631 38.007 61.681 ;
      RECT 35.477 61.585 38.053 61.635 ;
      RECT 35.523 61.539 38.099 61.589 ;
      RECT 35.569 61.493 38.145 61.543 ;
      RECT 35.615 61.447 38.191 61.497 ;
      RECT 35.661 61.401 38.237 61.451 ;
      RECT 35.707 61.355 38.283 61.405 ;
      RECT 35.753 61.309 38.329 61.359 ;
      RECT 35.799 61.263 38.375 61.313 ;
      RECT 35.845 61.217 38.421 61.267 ;
      RECT 35.891 61.171 38.467 61.221 ;
      RECT 35.937 61.125 38.513 61.175 ;
      RECT 35.983 61.079 38.559 61.129 ;
      RECT 36.029 61.033 38.605 61.083 ;
      RECT 36.075 60.987 38.651 61.037 ;
      RECT 36.121 60.941 38.697 60.991 ;
      RECT 36.167 60.895 38.743 60.945 ;
      RECT 36.213 60.849 38.789 60.899 ;
      RECT 36.259 60.803 38.835 60.853 ;
      RECT 36.305 60.757 38.881 60.807 ;
      RECT 36.351 60.711 38.927 60.761 ;
      RECT 36.397 60.665 38.973 60.715 ;
      RECT 36.443 60.619 39.019 60.669 ;
      RECT 36.489 60.573 39.065 60.623 ;
      RECT 36.535 60.527 39.111 60.577 ;
      RECT 36.581 60.481 39.157 60.531 ;
      RECT 36.627 60.435 39.203 60.485 ;
      RECT 36.673 60.389 39.249 60.439 ;
      RECT 36.719 60.343 39.295 60.393 ;
      RECT 36.765 60.297 39.341 60.347 ;
      RECT 36.811 60.251 39.387 60.301 ;
      RECT 36.857 60.205 39.433 60.255 ;
      RECT 36.903 60.159 39.479 60.209 ;
      RECT 36.949 60.113 39.525 60.163 ;
      RECT 36.995 60.067 39.571 60.117 ;
      RECT 37.041 60.021 39.617 60.071 ;
      RECT 37.087 59.975 39.663 60.025 ;
      RECT 37.133 59.929 39.709 59.979 ;
      RECT 37.179 59.883 39.755 59.933 ;
      RECT 37.225 59.837 39.801 59.887 ;
      RECT 37.271 59.791 39.847 59.841 ;
      RECT 37.317 59.745 39.893 59.795 ;
      RECT 37.363 59.699 39.939 59.749 ;
      RECT 37.409 59.653 39.985 59.703 ;
      RECT 37.455 59.607 40.031 59.657 ;
      RECT 37.501 59.561 40.077 59.611 ;
      RECT 37.547 59.515 40.123 59.565 ;
      RECT 37.593 59.469 40.169 59.519 ;
      RECT 37.639 59.423 40.215 59.473 ;
      RECT 37.685 59.377 40.261 59.427 ;
      RECT 37.731 59.331 40.307 59.381 ;
      RECT 37.777 59.285 40.353 59.335 ;
      RECT 37.823 59.239 40.399 59.289 ;
      RECT 37.869 59.193 40.445 59.243 ;
      RECT 37.915 59.147 40.491 59.197 ;
      RECT 37.961 59.101 40.537 59.151 ;
      RECT 38.007 59.055 40.583 59.105 ;
      RECT 38.053 59.009 40.629 59.059 ;
      RECT 38.099 58.963 40.675 59.013 ;
      RECT 38.145 58.917 40.721 58.967 ;
      RECT 38.191 58.871 40.767 58.921 ;
      RECT 38.237 58.825 40.813 58.875 ;
      RECT 38.283 58.779 40.859 58.829 ;
      RECT 38.329 58.733 40.905 58.783 ;
      RECT 38.375 58.687 40.951 58.737 ;
      RECT 38.421 58.641 40.997 58.691 ;
      RECT 38.467 58.595 41.043 58.645 ;
      RECT 38.513 58.549 41.089 58.599 ;
      RECT 38.559 58.503 41.135 58.553 ;
      RECT 38.605 58.457 41.181 58.507 ;
      RECT 38.651 58.411 41.227 58.461 ;
      RECT 38.697 58.365 41.273 58.415 ;
      RECT 38.743 58.319 41.319 58.369 ;
      RECT 38.789 58.273 41.365 58.323 ;
      RECT 38.835 58.227 41.411 58.277 ;
      RECT 38.881 58.181 41.457 58.231 ;
      RECT 38.927 58.135 41.503 58.185 ;
      RECT 38.973 58.089 41.549 58.139 ;
      RECT 39.019 58.043 41.595 58.093 ;
      RECT 39.065 57.997 41.641 58.047 ;
      RECT 39.111 57.951 41.687 58.001 ;
      RECT 39.157 57.905 41.733 57.955 ;
      RECT 39.203 57.859 41.779 57.909 ;
      RECT 39.249 57.813 41.825 57.863 ;
      RECT 39.295 57.767 41.871 57.817 ;
      RECT 39.341 57.721 41.917 57.771 ;
      RECT 39.387 57.675 41.963 57.725 ;
      RECT 39.433 57.629 42.009 57.679 ;
      RECT 39.479 57.583 42.055 57.633 ;
      RECT 39.525 57.537 42.101 57.587 ;
      RECT 39.571 57.491 42.147 57.541 ;
      RECT 39.617 57.445 42.193 57.495 ;
      RECT 39.663 57.399 42.239 57.449 ;
      RECT 39.709 57.353 42.285 57.403 ;
      RECT 39.755 57.307 42.325 57.36 ;
      RECT 39.801 57.261 42.371 57.317 ;
      RECT 39.847 57.215 42.417 57.271 ;
      RECT 39.893 57.169 42.463 57.225 ;
      RECT 39.939 57.123 42.509 57.179 ;
      RECT 39.985 57.077 42.555 57.133 ;
      RECT 40.031 57.031 42.601 57.087 ;
      RECT 40.077 56.985 42.647 57.041 ;
      RECT 40.123 56.939 42.693 56.995 ;
      RECT 40.169 56.893 42.739 56.949 ;
      RECT 40.215 56.847 42.785 56.903 ;
      RECT 40.261 56.801 42.831 56.857 ;
      RECT 40.307 56.755 42.877 56.811 ;
      RECT 40.353 56.709 42.923 56.765 ;
      RECT 40.399 56.663 42.969 56.719 ;
      RECT 40.445 56.617 43.015 56.673 ;
      RECT 40.491 56.571 43.061 56.627 ;
      RECT 40.537 56.525 43.107 56.581 ;
      RECT 40.583 56.479 43.153 56.535 ;
      RECT 40.629 56.433 43.199 56.489 ;
      RECT 40.675 56.387 43.245 56.443 ;
      RECT 40.721 56.341 43.291 56.397 ;
      RECT 40.767 56.295 43.337 56.351 ;
      RECT 40.813 56.249 43.383 56.305 ;
      RECT 40.859 56.203 43.429 56.259 ;
      RECT 40.905 56.157 43.475 56.213 ;
      RECT 40.951 56.111 43.521 56.167 ;
      RECT 40.997 56.065 43.567 56.121 ;
      RECT 41.043 56.019 43.613 56.075 ;
      RECT 41.089 55.973 43.659 56.029 ;
      RECT 41.135 55.927 43.705 55.983 ;
      RECT 41.181 55.881 43.751 55.937 ;
      RECT 41.227 55.835 43.797 55.891 ;
      RECT 41.273 55.789 43.843 55.845 ;
      RECT 41.319 55.743 43.889 55.799 ;
      RECT 41.365 55.697 43.935 55.753 ;
      RECT 41.411 55.651 43.981 55.707 ;
      RECT 41.457 55.605 44.027 55.661 ;
      RECT 41.503 55.559 44.073 55.615 ;
      RECT 41.549 55.513 44.119 55.569 ;
      RECT 41.595 55.467 44.165 55.523 ;
      RECT 41.641 55.421 44.211 55.477 ;
      RECT 41.687 55.375 44.257 55.431 ;
      RECT 41.733 55.329 44.303 55.385 ;
      RECT 41.779 55.283 44.349 55.339 ;
      RECT 41.825 55.237 44.395 55.293 ;
      RECT 41.871 55.191 44.441 55.247 ;
      RECT 41.917 55.145 44.487 55.201 ;
      RECT 41.963 55.099 44.533 55.155 ;
      RECT 42.009 55.053 44.579 55.109 ;
      RECT 42.055 55.007 44.625 55.063 ;
      RECT 42.101 54.961 44.671 55.017 ;
      RECT 42.147 54.915 44.717 54.971 ;
      RECT 42.193 54.869 44.763 54.925 ;
      RECT 42.239 54.823 44.809 54.879 ;
      RECT 42.285 54.777 44.855 54.833 ;
      RECT 42.331 54.731 44.901 54.787 ;
      RECT 42.377 54.685 44.947 54.741 ;
      RECT 42.423 54.639 44.993 54.695 ;
      RECT 42.469 54.593 45.039 54.649 ;
      RECT 42.515 54.547 45.085 54.603 ;
      RECT 42.561 54.501 45.131 54.557 ;
      RECT 42.607 54.455 45.177 54.511 ;
      RECT 42.653 54.409 45.223 54.465 ;
      RECT 42.699 54.363 45.269 54.419 ;
      RECT 42.745 54.317 45.315 54.373 ;
      RECT 42.791 54.271 45.361 54.327 ;
      RECT 42.837 54.225 45.407 54.281 ;
      RECT 42.883 54.179 45.453 54.235 ;
      RECT 42.929 54.133 45.499 54.189 ;
      RECT 42.975 54.087 45.545 54.143 ;
      RECT 43.021 54.041 45.591 54.097 ;
      RECT 43.067 53.995 45.637 54.051 ;
      RECT 43.113 53.949 45.683 54.005 ;
      RECT 43.159 53.903 45.729 53.959 ;
      RECT 43.205 53.857 45.775 53.913 ;
      RECT 43.251 53.811 45.821 53.867 ;
      RECT 43.297 53.765 45.867 53.821 ;
      RECT 43.343 53.719 45.913 53.775 ;
      RECT 43.389 53.673 45.959 53.729 ;
      RECT 43.435 53.627 46.005 53.683 ;
      RECT 43.481 53.581 46.051 53.637 ;
      RECT 43.527 53.535 46.097 53.591 ;
      RECT 43.573 53.489 46.143 53.545 ;
      RECT 43.619 53.443 46.189 53.499 ;
      RECT 43.665 53.397 46.235 53.453 ;
      RECT 43.711 53.351 46.281 53.407 ;
      RECT 43.757 53.305 46.327 53.361 ;
      RECT 43.803 53.259 46.373 53.315 ;
      RECT 43.849 53.213 46.419 53.269 ;
      RECT 43.895 53.167 46.465 53.223 ;
      RECT 43.941 53.121 46.511 53.177 ;
      RECT 43.987 53.075 46.557 53.131 ;
      RECT 44.033 53.029 46.603 53.085 ;
      RECT 44.079 52.983 46.649 53.039 ;
      RECT 44.125 52.937 46.695 52.993 ;
      RECT 44.171 52.891 46.741 52.947 ;
      RECT 44.217 52.845 46.787 52.901 ;
      RECT 44.263 52.799 46.833 52.855 ;
      RECT 44.309 52.753 46.879 52.809 ;
      RECT 44.355 52.707 46.925 52.763 ;
      RECT 44.401 52.661 46.971 52.717 ;
      RECT 44.447 52.615 47.017 52.671 ;
      RECT 44.493 52.569 47.063 52.625 ;
      RECT 44.539 52.523 47.109 52.579 ;
      RECT 44.585 52.477 47.155 52.533 ;
      RECT 44.631 52.431 47.201 52.487 ;
      RECT 44.677 52.385 47.247 52.441 ;
      RECT 44.723 52.339 47.293 52.395 ;
      RECT 44.769 52.293 47.339 52.349 ;
      RECT 44.815 52.247 47.385 52.303 ;
      RECT 44.861 52.201 47.431 52.257 ;
      RECT 44.907 52.155 47.477 52.211 ;
      RECT 44.953 52.109 47.523 52.165 ;
      RECT 44.999 52.063 47.569 52.119 ;
      RECT 45.045 52.017 47.615 52.073 ;
      RECT 45.091 51.971 47.661 52.027 ;
      RECT 45.137 51.925 47.707 51.981 ;
      RECT 45.183 51.879 47.753 51.935 ;
      RECT 45.229 51.833 47.799 51.889 ;
      RECT 45.275 51.787 47.845 51.843 ;
      RECT 45.321 51.741 47.891 51.797 ;
      RECT 45.367 51.695 47.937 51.751 ;
      RECT 45.413 51.649 47.983 51.705 ;
      RECT 45.459 51.603 48.029 51.659 ;
      RECT 45.505 51.557 48.075 51.613 ;
      RECT 45.551 51.511 48.121 51.567 ;
      RECT 45.597 51.465 48.167 51.521 ;
      RECT 45.643 51.419 48.213 51.475 ;
      RECT 45.689 51.373 48.259 51.429 ;
      RECT 45.735 51.327 48.305 51.383 ;
      RECT 45.781 51.281 48.351 51.337 ;
      RECT 45.827 51.235 48.397 51.291 ;
      RECT 45.873 51.189 48.443 51.245 ;
      RECT 45.919 51.143 48.489 51.199 ;
      RECT 45.965 51.097 48.535 51.153 ;
      RECT 46.011 51.051 48.581 51.107 ;
      RECT 46.057 51.005 48.627 51.061 ;
      RECT 46.103 50.959 48.673 51.015 ;
      RECT 46.149 50.913 48.719 50.969 ;
      RECT 46.195 50.867 48.765 50.923 ;
      RECT 46.241 50.821 48.811 50.877 ;
      RECT 46.287 50.775 48.857 50.831 ;
      RECT 46.333 50.729 48.903 50.785 ;
      RECT 46.379 50.683 48.949 50.739 ;
      RECT 46.425 50.637 48.995 50.693 ;
      RECT 46.471 50.591 49.041 50.647 ;
      RECT 46.517 50.545 49.087 50.601 ;
      RECT 46.563 50.499 49.133 50.555 ;
      RECT 46.609 50.453 49.179 50.509 ;
      RECT 46.655 50.407 49.225 50.463 ;
      RECT 46.701 50.361 49.271 50.417 ;
      RECT 46.747 50.315 49.317 50.371 ;
      RECT 46.793 50.269 49.363 50.325 ;
      RECT 46.839 50.223 49.409 50.279 ;
      RECT 46.885 50.177 49.455 50.233 ;
      RECT 46.931 50.131 49.501 50.187 ;
      RECT 46.977 50.085 49.547 50.141 ;
      RECT 47.023 50.039 49.593 50.095 ;
      RECT 47.069 49.993 49.639 50.049 ;
      RECT 47.115 49.947 49.685 50.003 ;
      RECT 47.161 49.901 49.731 49.957 ;
      RECT 47.207 49.855 49.777 49.911 ;
      RECT 47.253 49.809 49.823 49.865 ;
      RECT 47.299 49.763 49.869 49.819 ;
      RECT 47.345 49.717 49.915 49.773 ;
      RECT 47.391 49.671 49.961 49.727 ;
      RECT 47.437 49.625 50.007 49.681 ;
      RECT 47.483 49.579 50.053 49.635 ;
      RECT 47.529 49.533 50.099 49.589 ;
      RECT 47.575 49.487 50.145 49.543 ;
      RECT 47.621 49.441 50.191 49.497 ;
      RECT 47.667 49.395 50.237 49.451 ;
      RECT 47.713 49.349 50.283 49.405 ;
      RECT 47.759 49.303 50.329 49.359 ;
      RECT 47.805 49.257 50.375 49.313 ;
      RECT 47.851 49.211 50.421 49.267 ;
      RECT 47.897 49.165 50.467 49.221 ;
      RECT 47.943 49.119 50.513 49.175 ;
      RECT 47.989 49.073 50.559 49.129 ;
      RECT 48.035 49.027 50.605 49.083 ;
      RECT 48.081 48.981 50.651 49.037 ;
      RECT 48.127 48.935 50.697 48.991 ;
      RECT 48.173 48.889 50.743 48.945 ;
      RECT 48.219 48.843 50.789 48.899 ;
      RECT 48.265 48.797 50.835 48.853 ;
      RECT 48.311 48.751 50.881 48.807 ;
      RECT 48.357 48.705 50.927 48.761 ;
      RECT 48.403 48.659 50.973 48.715 ;
      RECT 48.449 48.613 51.019 48.669 ;
      RECT 48.495 48.567 51.065 48.623 ;
      RECT 48.541 48.521 51.111 48.577 ;
      RECT 48.587 48.475 51.157 48.531 ;
      RECT 48.633 48.429 51.203 48.485 ;
      RECT 48.679 48.383 51.249 48.439 ;
      RECT 48.725 48.337 51.295 48.393 ;
      RECT 48.771 48.291 51.341 48.347 ;
      RECT 48.817 48.245 51.387 48.301 ;
      RECT 48.863 48.199 51.433 48.255 ;
      RECT 48.909 48.153 51.479 48.209 ;
      RECT 48.955 48.107 51.525 48.163 ;
      RECT 49.001 48.061 51.571 48.117 ;
      RECT 49.047 48.015 51.617 48.071 ;
      RECT 49.093 47.969 51.663 48.025 ;
      RECT 49.139 47.923 51.709 47.979 ;
      RECT 49.185 47.877 51.755 47.933 ;
      RECT 49.231 47.831 51.801 47.887 ;
      RECT 49.277 47.785 51.847 47.841 ;
      RECT 49.323 47.739 51.893 47.795 ;
      RECT 49.369 47.693 51.939 47.749 ;
      RECT 49.415 47.647 51.985 47.703 ;
      RECT 49.461 47.601 52.031 47.657 ;
      RECT 49.507 47.555 52.077 47.611 ;
      RECT 49.553 47.509 52.123 47.565 ;
      RECT 49.599 47.463 52.169 47.519 ;
      RECT 49.645 47.417 52.215 47.473 ;
      RECT 49.691 47.371 52.261 47.427 ;
      RECT 49.737 47.325 52.307 47.381 ;
      RECT 49.783 47.279 52.353 47.335 ;
      RECT 49.829 47.233 52.399 47.289 ;
      RECT 49.875 47.187 52.445 47.243 ;
      RECT 49.921 47.141 52.491 47.197 ;
      RECT 49.967 47.095 52.537 47.151 ;
      RECT 50.013 47.049 52.583 47.105 ;
      RECT 50.059 47.003 52.629 47.059 ;
      RECT 50.105 46.957 52.675 47.013 ;
      RECT 50.151 46.911 52.721 46.967 ;
      RECT 50.197 46.865 52.767 46.921 ;
      RECT 50.243 46.819 52.813 46.875 ;
      RECT 50.289 46.773 52.859 46.829 ;
      RECT 50.335 46.727 52.905 46.783 ;
      RECT 50.381 46.681 52.951 46.737 ;
      RECT 50.427 46.635 52.997 46.691 ;
      RECT 50.473 46.589 53.043 46.645 ;
      RECT 50.519 46.543 53.089 46.599 ;
      RECT 50.565 46.497 53.135 46.553 ;
      RECT 50.611 46.451 53.181 46.507 ;
      RECT 50.657 46.405 53.227 46.461 ;
      RECT 50.703 46.359 53.273 46.415 ;
      RECT 50.749 46.313 53.319 46.369 ;
      RECT 50.795 46.267 53.365 46.323 ;
      RECT 50.841 46.221 53.411 46.277 ;
      RECT 50.887 46.175 53.457 46.231 ;
      RECT 50.933 46.129 53.503 46.185 ;
      RECT 50.979 46.083 53.549 46.139 ;
      RECT 51.025 46.037 53.595 46.093 ;
      RECT 51.071 45.991 53.641 46.047 ;
      RECT 51.117 45.945 53.687 46.001 ;
      RECT 51.163 45.899 53.733 45.955 ;
      RECT 51.209 45.853 53.779 45.909 ;
      RECT 51.255 45.807 53.825 45.863 ;
      RECT 51.301 45.761 53.871 45.817 ;
      RECT 51.347 45.715 53.917 45.771 ;
      RECT 51.393 45.669 53.963 45.725 ;
      RECT 51.439 45.623 54.009 45.679 ;
      RECT 51.485 45.577 54.055 45.633 ;
      RECT 51.531 45.531 54.101 45.587 ;
      RECT 51.577 45.485 54.147 45.541 ;
      RECT 51.623 45.439 54.193 45.495 ;
      RECT 51.669 45.393 54.239 45.449 ;
      RECT 51.715 45.347 54.285 45.403 ;
      RECT 51.761 45.301 54.331 45.357 ;
      RECT 51.807 45.255 54.377 45.311 ;
      RECT 51.853 45.209 54.423 45.265 ;
      RECT 51.899 45.163 54.469 45.219 ;
      RECT 51.945 45.117 54.515 45.173 ;
      RECT 51.991 45.071 54.561 45.127 ;
      RECT 52.037 45.025 54.607 45.081 ;
      RECT 52.083 44.979 54.653 45.035 ;
      RECT 52.129 44.933 54.699 44.989 ;
      RECT 52.175 44.887 54.745 44.943 ;
      RECT 52.221 44.841 54.791 44.897 ;
      RECT 52.267 44.795 54.837 44.851 ;
      RECT 52.313 44.749 54.883 44.805 ;
      RECT 52.359 44.703 54.929 44.759 ;
      RECT 52.405 44.657 54.975 44.713 ;
      RECT 52.451 44.611 55.021 44.667 ;
      RECT 52.497 44.565 55.067 44.621 ;
      RECT 52.543 44.519 55.113 44.575 ;
      RECT 52.589 44.473 55.159 44.529 ;
      RECT 52.635 44.427 55.205 44.483 ;
      RECT 52.681 44.381 55.251 44.437 ;
      RECT 52.727 44.335 55.297 44.391 ;
      RECT 52.773 44.289 55.343 44.345 ;
      RECT 52.819 44.243 55.389 44.299 ;
      RECT 52.865 44.197 55.435 44.253 ;
      RECT 52.911 44.151 55.481 44.207 ;
      RECT 52.957 44.105 55.527 44.161 ;
      RECT 53.003 44.059 55.573 44.115 ;
      RECT 53.049 44.013 55.619 44.069 ;
      RECT 53.095 43.967 55.665 44.023 ;
      RECT 53.141 43.921 55.711 43.977 ;
      RECT 53.187 43.875 55.757 43.931 ;
      RECT 53.233 43.829 55.803 43.885 ;
      RECT 53.279 43.783 55.849 43.839 ;
      RECT 53.325 43.737 55.895 43.793 ;
      RECT 53.371 43.691 55.941 43.747 ;
      RECT 53.417 43.645 55.987 43.701 ;
      RECT 53.463 43.599 56.033 43.655 ;
      RECT 53.509 43.553 56.079 43.609 ;
      RECT 53.555 43.507 56.125 43.563 ;
      RECT 53.601 43.461 56.171 43.517 ;
      RECT 53.647 43.415 56.217 43.471 ;
      RECT 53.693 43.369 56.263 43.425 ;
      RECT 53.739 43.323 56.309 43.379 ;
      RECT 53.785 43.277 56.355 43.333 ;
      RECT 53.831 43.231 56.401 43.287 ;
      RECT 53.877 43.185 56.447 43.241 ;
      RECT 53.923 43.139 56.493 43.195 ;
      RECT 53.969 43.093 56.539 43.149 ;
      RECT 54.015 43.047 56.585 43.103 ;
      RECT 54.061 43.001 56.631 43.057 ;
      RECT 54.107 42.955 56.677 43.011 ;
      RECT 54.153 42.909 56.723 42.965 ;
      RECT 54.199 42.863 56.769 42.919 ;
      RECT 54.245 42.817 56.815 42.873 ;
      RECT 54.291 42.771 56.861 42.827 ;
      RECT 54.337 42.725 56.907 42.781 ;
      RECT 54.383 42.679 56.953 42.735 ;
      RECT 54.429 42.633 56.999 42.689 ;
      RECT 54.475 42.587 57.045 42.643 ;
      RECT 54.521 42.541 57.091 42.597 ;
      RECT 54.567 42.495 57.137 42.551 ;
      RECT 54.613 42.449 57.183 42.505 ;
      RECT 54.659 42.403 57.229 42.459 ;
      RECT 54.705 42.357 57.275 42.413 ;
      RECT 54.751 42.311 57.321 42.367 ;
      RECT 54.797 42.265 57.367 42.321 ;
      RECT 54.843 42.219 57.413 42.275 ;
      RECT 54.889 42.173 57.459 42.229 ;
      RECT 54.935 42.127 57.505 42.183 ;
      RECT 54.981 42.081 57.551 42.137 ;
      RECT 55.027 42.035 57.597 42.091 ;
      RECT 55.073 41.989 57.643 42.045 ;
      RECT 55.119 41.943 57.689 41.999 ;
      RECT 55.165 41.897 57.735 41.953 ;
      RECT 55.211 41.851 57.781 41.907 ;
      RECT 55.257 41.805 57.827 41.861 ;
      RECT 55.303 41.759 57.873 41.815 ;
      RECT 55.349 41.713 57.919 41.769 ;
      RECT 55.395 41.667 57.965 41.723 ;
      RECT 55.441 41.621 58.011 41.677 ;
      RECT 55.487 41.575 58.057 41.631 ;
      RECT 55.533 41.529 58.103 41.585 ;
      RECT 55.579 41.483 58.149 41.539 ;
      RECT 55.625 41.437 58.195 41.493 ;
      RECT 55.671 41.391 58.241 41.447 ;
      RECT 55.717 41.345 58.287 41.401 ;
      RECT 55.763 41.299 58.333 41.355 ;
      RECT 55.809 41.253 58.379 41.309 ;
      RECT 55.855 41.207 58.425 41.263 ;
      RECT 55.901 41.161 58.471 41.217 ;
      RECT 55.947 41.115 58.517 41.171 ;
      RECT 55.993 41.069 58.563 41.125 ;
      RECT 56.039 41.023 58.609 41.079 ;
      RECT 56.085 40.977 58.655 41.033 ;
      RECT 56.131 40.931 58.701 40.987 ;
      RECT 56.177 40.885 58.747 40.941 ;
      RECT 56.223 40.839 58.793 40.895 ;
      RECT 56.269 40.793 58.839 40.849 ;
      RECT 56.315 40.747 58.885 40.803 ;
      RECT 56.361 40.701 58.931 40.757 ;
      RECT 56.407 40.655 58.977 40.711 ;
      RECT 56.453 40.609 59.023 40.665 ;
      RECT 56.499 40.563 59.069 40.619 ;
      RECT 56.545 40.517 59.115 40.573 ;
      RECT 56.591 40.471 59.161 40.527 ;
      RECT 56.637 40.425 59.207 40.481 ;
      RECT 56.683 40.379 59.253 40.435 ;
      RECT 56.729 40.333 59.299 40.389 ;
      RECT 56.775 40.287 59.345 40.343 ;
      RECT 56.821 40.241 59.391 40.297 ;
      RECT 56.867 40.195 59.437 40.251 ;
      RECT 56.913 40.149 59.483 40.205 ;
      RECT 56.959 40.103 59.529 40.159 ;
      RECT 57.005 40.057 59.575 40.113 ;
      RECT 57.051 40.011 59.621 40.067 ;
      RECT 57.097 39.965 59.667 40.021 ;
      RECT 57.143 39.919 59.713 39.975 ;
      RECT 57.189 39.873 59.759 39.929 ;
      RECT 57.235 39.827 59.805 39.883 ;
      RECT 57.281 39.781 59.851 39.837 ;
      RECT 57.327 39.735 59.897 39.791 ;
      RECT 57.373 39.689 59.943 39.745 ;
      RECT 57.419 39.643 59.989 39.699 ;
      RECT 57.465 39.597 60.035 39.653 ;
      RECT 57.511 39.551 60.081 39.607 ;
      RECT 57.557 39.505 60.127 39.561 ;
      RECT 57.603 39.459 60.173 39.515 ;
      RECT 57.649 39.413 60.219 39.469 ;
      RECT 57.695 39.367 60.265 39.423 ;
      RECT 57.741 39.321 60.311 39.377 ;
      RECT 57.787 39.275 60.357 39.331 ;
      RECT 57.833 39.229 60.403 39.285 ;
      RECT 57.879 39.183 60.449 39.239 ;
      RECT 57.925 39.137 60.495 39.193 ;
      RECT 57.971 39.091 60.541 39.147 ;
      RECT 58.017 39.045 60.587 39.101 ;
      RECT 58.063 38.999 60.633 39.055 ;
      RECT 58.109 38.953 60.679 39.009 ;
      RECT 58.155 38.907 60.725 38.963 ;
      RECT 58.201 38.861 60.771 38.917 ;
      RECT 58.247 38.815 60.817 38.871 ;
      RECT 58.293 38.769 60.863 38.825 ;
      RECT 58.339 38.723 60.909 38.779 ;
      RECT 58.385 38.677 60.955 38.733 ;
      RECT 58.431 38.631 61.001 38.687 ;
      RECT 58.477 38.585 61.047 38.641 ;
      RECT 58.523 38.539 61.093 38.595 ;
      RECT 58.569 38.493 61.139 38.549 ;
      RECT 58.615 38.447 61.185 38.503 ;
      RECT 58.661 38.401 61.231 38.457 ;
      RECT 58.707 38.355 61.277 38.411 ;
      RECT 58.753 38.309 61.323 38.365 ;
      RECT 58.799 38.263 61.369 38.319 ;
      RECT 58.845 38.217 61.415 38.273 ;
      RECT 58.891 38.171 61.461 38.227 ;
      RECT 58.937 38.125 61.507 38.181 ;
      RECT 58.983 38.079 61.553 38.135 ;
      RECT 59.029 38.033 61.599 38.089 ;
      RECT 59.075 37.987 61.645 38.043 ;
      RECT 59.121 37.941 61.691 37.997 ;
      RECT 59.167 37.895 61.737 37.951 ;
      RECT 59.213 37.849 61.783 37.905 ;
      RECT 59.259 37.803 61.829 37.859 ;
      RECT 59.305 37.757 61.875 37.813 ;
      RECT 59.351 37.711 61.921 37.767 ;
      RECT 59.397 37.665 61.967 37.721 ;
      RECT 59.443 37.619 62.013 37.675 ;
      RECT 59.489 37.573 62.059 37.629 ;
      RECT 59.535 37.527 62.105 37.583 ;
      RECT 59.581 37.481 62.151 37.537 ;
      RECT 59.627 37.435 62.197 37.491 ;
      RECT 59.673 37.389 62.243 37.445 ;
      RECT 59.719 37.343 62.289 37.399 ;
      RECT 59.765 37.297 62.335 37.353 ;
      RECT 59.811 37.251 62.381 37.307 ;
      RECT 59.857 37.205 62.427 37.261 ;
      RECT 59.903 37.159 62.473 37.215 ;
      RECT 59.949 37.113 62.519 37.169 ;
      RECT 59.995 37.067 62.565 37.123 ;
      RECT 60.041 37.021 62.611 37.077 ;
      RECT 60.087 36.975 62.657 37.031 ;
      RECT 60.133 36.929 62.703 36.985 ;
      RECT 60.179 36.883 62.749 36.939 ;
      RECT 60.225 36.837 62.795 36.893 ;
      RECT 60.271 36.791 62.841 36.847 ;
      RECT 60.317 36.745 62.887 36.801 ;
      RECT 60.363 36.699 62.933 36.755 ;
      RECT 60.409 36.653 62.979 36.709 ;
      RECT 62.939 34.146 62.979 36.709 ;
      RECT 60.455 36.607 63.025 36.663 ;
      RECT 62.94 34.122 63.025 36.663 ;
      RECT 60.501 36.561 63.071 36.617 ;
      RECT 62.986 34.076 63.071 36.617 ;
      RECT 60.547 36.515 63.117 36.571 ;
      RECT 63.032 34.03 63.117 36.571 ;
      RECT 60.593 36.469 63.163 36.525 ;
      RECT 63.078 33.984 63.163 36.525 ;
      RECT 60.639 36.423 63.209 36.479 ;
      RECT 63.124 33.938 63.209 36.479 ;
      RECT 60.685 36.377 63.255 36.433 ;
      RECT 63.17 33.892 63.255 36.433 ;
      RECT 60.731 36.331 63.301 36.387 ;
      RECT 63.216 33.846 63.301 36.387 ;
      RECT 60.777 36.285 63.347 36.341 ;
      RECT 63.262 33.8 63.347 36.341 ;
      RECT 60.823 36.239 63.393 36.295 ;
      RECT 63.308 33.754 63.393 36.295 ;
      RECT 60.869 36.193 63.439 36.249 ;
      RECT 63.354 33.708 63.439 36.249 ;
      RECT 60.915 36.147 63.485 36.203 ;
      RECT 63.4 33.662 63.485 36.203 ;
      RECT 60.961 36.101 63.531 36.157 ;
      RECT 63.446 33.616 63.531 36.157 ;
      RECT 61.007 36.055 63.577 36.111 ;
      RECT 63.492 33.57 63.577 36.111 ;
      RECT 61.053 36.009 63.623 36.065 ;
      RECT 63.538 33.524 63.623 36.065 ;
      RECT 61.099 35.963 63.669 36.019 ;
      RECT 63.584 33.478 63.669 36.019 ;
      RECT 61.145 35.917 63.715 35.973 ;
      RECT 63.63 33.432 63.715 35.973 ;
      RECT 61.191 35.871 63.761 35.927 ;
      RECT 63.676 33.386 63.761 35.927 ;
      RECT 61.237 35.825 63.807 35.881 ;
      RECT 63.722 33.34 63.807 35.881 ;
      RECT 61.283 35.779 63.853 35.835 ;
      RECT 63.768 33.294 63.853 35.835 ;
      RECT 61.329 35.733 63.899 35.789 ;
      RECT 63.814 33.248 63.899 35.789 ;
      RECT 61.375 35.687 63.945 35.743 ;
      RECT 63.86 33.202 63.945 35.743 ;
      RECT 61.421 35.641 63.991 35.697 ;
      RECT 63.906 33.156 63.991 35.697 ;
      RECT 61.467 35.595 64.037 35.651 ;
      RECT 63.952 33.11 64.037 35.651 ;
      RECT 61.513 35.549 64.083 35.605 ;
      RECT 63.998 33.064 64.083 35.605 ;
      RECT 61.559 35.503 64.129 35.559 ;
      RECT 64.044 33.018 64.129 35.559 ;
      RECT 61.605 35.457 64.175 35.513 ;
      RECT 64.09 32.972 64.175 35.513 ;
      RECT 61.651 35.411 64.221 35.467 ;
      RECT 64.136 32.926 64.221 35.467 ;
      RECT 61.697 35.365 64.267 35.421 ;
      RECT 64.182 32.88 64.267 35.421 ;
      RECT 61.743 35.319 64.313 35.375 ;
      RECT 64.228 32.834 64.313 35.375 ;
      RECT 61.789 35.273 64.359 35.329 ;
      RECT 64.274 32.788 64.359 35.329 ;
      RECT 61.835 35.227 64.405 35.283 ;
      RECT 64.32 32.742 64.405 35.283 ;
      RECT 61.881 35.181 64.451 35.237 ;
      RECT 64.366 32.696 64.451 35.237 ;
      RECT 61.927 35.135 64.497 35.191 ;
      RECT 64.412 32.65 64.497 35.191 ;
      RECT 61.973 35.089 64.543 35.145 ;
      RECT 64.458 32.604 64.543 35.145 ;
      RECT 62.019 35.043 64.589 35.099 ;
      RECT 64.504 32.558 64.589 35.099 ;
      RECT 62.065 34.997 64.635 35.053 ;
      RECT 64.55 32.512 64.635 35.053 ;
      RECT 62.111 34.951 64.681 35.007 ;
      RECT 64.596 32.466 64.681 35.007 ;
      RECT 62.157 34.905 64.727 34.961 ;
      RECT 64.642 32.42 64.727 34.961 ;
      RECT 62.203 34.859 64.773 34.915 ;
      RECT 64.688 32.374 64.773 34.915 ;
      RECT 62.249 34.813 64.819 34.869 ;
      RECT 64.734 32.328 64.819 34.869 ;
      RECT 62.295 34.767 64.865 34.823 ;
      RECT 64.78 32.282 64.865 34.823 ;
      RECT 62.341 34.721 64.911 34.777 ;
      RECT 64.826 32.236 64.911 34.777 ;
      RECT 62.387 34.675 64.957 34.731 ;
      RECT 64.872 32.19 64.957 34.731 ;
      RECT 62.433 34.629 65.003 34.685 ;
      RECT 64.918 32.144 65.003 34.685 ;
      RECT 62.479 34.583 65.049 34.639 ;
      RECT 64.964 32.098 65.049 34.639 ;
      RECT 62.525 34.537 65.095 34.593 ;
      RECT 65.01 32.052 65.095 34.593 ;
      RECT 62.571 34.491 65.141 34.547 ;
      RECT 65.056 32.006 65.141 34.547 ;
      RECT 62.617 34.445 65.187 34.501 ;
      RECT 65.102 31.96 65.187 34.501 ;
      RECT 62.663 34.399 65.233 34.455 ;
      RECT 65.148 31.914 65.233 34.455 ;
      RECT 62.709 34.353 65.279 34.409 ;
      RECT 65.194 31.868 65.279 34.409 ;
      RECT 62.755 34.307 65.325 34.363 ;
      RECT 65.24 31.822 65.325 34.363 ;
      RECT 62.801 34.261 65.371 34.317 ;
      RECT 65.286 31.776 65.371 34.317 ;
      RECT 62.847 34.215 65.417 34.271 ;
      RECT 65.332 31.73 65.417 34.271 ;
      RECT 62.893 34.169 65.463 34.225 ;
      RECT 65.378 31.684 65.463 34.225 ;
      RECT 65.424 31.638 65.509 34.179 ;
      RECT 65.47 31.592 65.555 34.133 ;
      RECT 65.516 31.546 65.601 34.087 ;
      RECT 65.562 31.5 65.647 34.041 ;
      RECT 65.608 31.454 65.693 33.995 ;
      RECT 65.654 31.408 65.739 33.949 ;
      RECT 65.7 31.362 65.785 33.903 ;
      RECT 65.746 31.316 65.831 33.857 ;
      RECT 65.792 31.27 65.877 33.811 ;
      RECT 65.838 31.224 65.923 33.765 ;
      RECT 65.884 31.178 65.969 33.719 ;
      RECT 65.93 31.132 66.015 33.673 ;
      RECT 65.976 31.086 66.061 33.627 ;
      RECT 66.022 31.04 66.107 33.581 ;
      RECT 66.068 30.994 66.153 33.535 ;
      RECT 66.114 30.948 66.199 33.489 ;
      RECT 66.16 30.902 66.245 33.443 ;
      RECT 66.206 30.856 66.291 33.397 ;
      RECT 66.252 30.81 66.337 33.351 ;
      RECT 66.298 30.764 66.383 33.305 ;
      RECT 66.344 30.718 66.429 33.259 ;
      RECT 66.39 30.672 66.475 33.213 ;
      RECT 66.436 30.626 66.521 33.167 ;
      RECT 66.482 30.58 66.567 33.121 ;
      RECT 66.528 30.534 66.613 33.075 ;
      RECT 66.574 30.488 66.659 33.029 ;
      RECT 66.62 30.442 66.705 32.983 ;
      RECT 66.666 30.396 66.751 32.937 ;
      RECT 66.712 30.35 66.797 32.891 ;
      RECT 66.758 30.304 66.843 32.845 ;
      RECT 66.804 30.258 66.889 32.799 ;
      RECT 66.85 30.212 66.935 32.753 ;
      RECT 66.896 30.166 66.981 32.707 ;
      RECT 66.942 30.12 67.027 32.661 ;
      RECT 66.988 30.074 67.073 32.615 ;
      RECT 67.034 30.028 67.119 32.569 ;
      RECT 67.08 29.982 67.165 32.523 ;
      RECT 67.126 29.936 67.211 32.477 ;
      RECT 67.172 29.89 67.257 32.431 ;
      RECT 67.218 29.844 67.303 32.385 ;
      RECT 67.264 29.798 67.349 32.339 ;
      RECT 67.31 29.752 67.395 32.293 ;
      RECT 67.356 29.706 67.441 32.247 ;
      RECT 67.402 29.66 67.487 32.201 ;
      RECT 67.448 29.614 67.533 32.155 ;
      RECT 67.494 29.568 67.579 32.109 ;
      RECT 67.54 29.522 67.625 32.063 ;
      RECT 67.586 29.476 67.671 32.017 ;
      RECT 67.632 29.43 67.717 31.971 ;
      RECT 67.678 29.384 67.763 31.925 ;
      RECT 67.724 29.338 67.809 31.879 ;
      RECT 67.77 29.292 67.855 31.833 ;
      RECT 67.816 29.246 67.901 31.787 ;
      RECT 67.862 29.199 67.947 31.741 ;
      RECT 67.908 29.175 67.993 31.695 ;
      RECT 67.908 29.175 68.039 31.649 ;
      RECT 67.908 29.175 68.085 31.603 ;
      RECT 67.908 29.175 68.131 31.557 ;
      RECT 67.908 29.175 68.177 31.511 ;
      RECT 67.908 29.175 68.223 31.465 ;
      RECT 67.908 29.175 68.269 31.419 ;
      RECT 67.908 29.175 68.315 31.373 ;
      RECT 67.908 29.175 68.361 31.327 ;
      RECT 67.908 29.175 68.407 31.281 ;
      RECT 67.908 29.175 68.453 31.235 ;
      RECT 67.908 29.175 68.499 31.189 ;
      RECT 67.908 29.175 68.545 31.143 ;
      RECT 67.908 29.175 68.591 31.097 ;
      RECT 67.908 29.175 68.637 31.051 ;
      RECT 67.908 29.175 68.683 31.005 ;
      RECT 67.908 29.175 68.729 30.959 ;
      RECT 67.908 29.175 68.775 30.913 ;
      RECT 67.908 29.175 68.821 30.867 ;
      RECT 67.908 29.175 68.867 30.821 ;
      RECT 67.908 29.175 68.913 30.775 ;
      RECT 67.908 29.175 68.959 30.729 ;
      RECT 67.908 29.175 69.005 30.683 ;
      RECT 67.908 29.175 69.051 30.637 ;
      RECT 67.908 29.175 69.097 30.591 ;
      RECT 67.908 29.175 69.143 30.545 ;
      RECT 67.908 29.175 69.189 30.499 ;
      RECT 67.908 29.175 69.235 30.453 ;
      RECT 67.908 29.175 69.281 30.407 ;
      RECT 67.908 29.175 69.327 30.361 ;
      RECT 66.758 30.304 69.34 30.331 ;
      RECT 67.908 29.175 110 30.325 ;
      RECT 42.675 74.637 43.825 110 ;
      RECT 42.675 74.637 43.871 76.067 ;
      RECT 42.675 74.637 43.917 76.021 ;
      RECT 42.675 74.637 43.963 75.975 ;
      RECT 42.675 74.637 44.009 75.929 ;
      RECT 42.675 74.637 44.055 75.883 ;
      RECT 42.675 74.637 44.101 75.837 ;
      RECT 42.675 74.637 44.147 75.791 ;
      RECT 42.675 74.637 44.193 75.745 ;
      RECT 42.675 74.637 44.239 75.699 ;
      RECT 42.675 74.637 44.285 75.653 ;
      RECT 42.675 74.637 44.331 75.607 ;
      RECT 42.675 74.637 44.377 75.561 ;
      RECT 42.675 74.637 44.423 75.515 ;
      RECT 42.675 74.637 44.469 75.469 ;
      RECT 42.675 74.637 44.515 75.423 ;
      RECT 42.675 74.637 44.561 75.377 ;
      RECT 42.675 74.637 44.607 75.331 ;
      RECT 42.675 74.637 44.653 75.285 ;
      RECT 42.675 74.637 44.699 75.239 ;
      RECT 42.675 74.637 44.745 75.193 ;
      RECT 42.675 74.637 44.791 75.147 ;
      RECT 42.675 74.637 44.837 75.101 ;
      RECT 42.675 74.637 44.883 75.055 ;
      RECT 42.675 74.637 44.929 75.009 ;
      RECT 42.675 74.637 44.975 74.963 ;
      RECT 42.675 74.637 45.021 74.917 ;
      RECT 42.675 74.637 45.067 74.871 ;
      RECT 42.675 74.637 45.113 74.825 ;
      RECT 42.675 74.637 45.159 74.779 ;
      RECT 42.675 74.637 45.205 74.733 ;
      RECT 42.675 74.637 45.251 74.687 ;
      RECT 42.721 74.591 45.297 74.641 ;
      RECT 42.767 74.545 45.343 74.595 ;
      RECT 42.813 74.499 45.389 74.549 ;
      RECT 42.859 74.453 45.435 74.503 ;
      RECT 42.905 74.407 45.481 74.457 ;
      RECT 42.951 74.361 45.527 74.411 ;
      RECT 42.997 74.315 45.573 74.365 ;
      RECT 43.043 74.269 45.619 74.319 ;
      RECT 43.089 74.223 45.665 74.273 ;
      RECT 43.135 74.177 45.711 74.227 ;
      RECT 43.181 74.131 45.757 74.181 ;
      RECT 43.227 74.085 45.803 74.135 ;
      RECT 43.273 74.039 45.849 74.089 ;
      RECT 43.319 73.993 45.895 74.043 ;
      RECT 43.365 73.947 45.941 73.997 ;
      RECT 43.411 73.901 45.987 73.951 ;
      RECT 43.457 73.855 46.033 73.905 ;
      RECT 43.503 73.809 46.079 73.859 ;
      RECT 43.549 73.763 46.125 73.813 ;
      RECT 43.595 73.717 46.171 73.767 ;
      RECT 43.641 73.671 46.217 73.721 ;
      RECT 43.687 73.625 46.263 73.675 ;
      RECT 43.733 73.579 46.309 73.629 ;
      RECT 43.779 73.533 46.355 73.583 ;
      RECT 43.825 73.487 46.401 73.537 ;
      RECT 43.871 73.441 46.447 73.491 ;
      RECT 43.917 73.395 46.493 73.445 ;
      RECT 43.963 73.349 46.539 73.399 ;
      RECT 44.009 73.303 46.585 73.353 ;
      RECT 44.055 73.257 46.631 73.307 ;
      RECT 44.101 73.211 46.677 73.261 ;
      RECT 44.147 73.165 46.723 73.215 ;
      RECT 44.193 73.119 46.769 73.169 ;
      RECT 44.239 73.073 46.815 73.123 ;
      RECT 44.285 73.027 46.861 73.077 ;
      RECT 44.331 72.981 46.907 73.031 ;
      RECT 44.377 72.935 46.953 72.985 ;
      RECT 44.423 72.889 46.999 72.939 ;
      RECT 44.469 72.843 47.045 72.893 ;
      RECT 44.515 72.797 47.091 72.847 ;
      RECT 44.561 72.751 47.137 72.801 ;
      RECT 44.607 72.705 47.183 72.755 ;
      RECT 44.653 72.659 47.229 72.709 ;
      RECT 44.699 72.613 47.275 72.663 ;
      RECT 44.745 72.567 47.321 72.617 ;
      RECT 44.791 72.521 47.367 72.571 ;
      RECT 44.837 72.475 47.413 72.525 ;
      RECT 44.883 72.429 47.459 72.479 ;
      RECT 44.929 72.383 47.505 72.433 ;
      RECT 44.975 72.337 47.551 72.387 ;
      RECT 45.021 72.291 47.597 72.341 ;
      RECT 45.067 72.245 47.643 72.295 ;
      RECT 45.113 72.199 47.689 72.249 ;
      RECT 45.159 72.153 47.735 72.203 ;
      RECT 45.205 72.107 47.781 72.157 ;
      RECT 45.251 72.061 47.827 72.111 ;
      RECT 45.297 72.015 47.873 72.065 ;
      RECT 45.343 71.969 47.919 72.019 ;
      RECT 45.389 71.923 47.965 71.973 ;
      RECT 45.435 71.877 48.011 71.927 ;
      RECT 45.481 71.831 48.057 71.881 ;
      RECT 45.527 71.785 48.103 71.835 ;
      RECT 45.573 71.739 48.149 71.789 ;
      RECT 45.619 71.693 48.195 71.743 ;
      RECT 45.665 71.647 48.241 71.697 ;
      RECT 45.711 71.601 48.287 71.651 ;
      RECT 45.757 71.555 48.333 71.605 ;
      RECT 45.803 71.509 48.379 71.559 ;
      RECT 45.849 71.463 48.425 71.513 ;
      RECT 45.895 71.417 48.471 71.467 ;
      RECT 45.941 71.371 48.517 71.421 ;
      RECT 45.987 71.325 48.563 71.375 ;
      RECT 46.033 71.279 48.609 71.329 ;
      RECT 46.079 71.233 48.655 71.283 ;
      RECT 46.125 71.187 48.701 71.237 ;
      RECT 46.171 71.141 48.747 71.191 ;
      RECT 46.217 71.095 48.793 71.145 ;
      RECT 46.263 71.049 48.839 71.099 ;
      RECT 46.309 71.003 48.885 71.053 ;
      RECT 46.355 70.957 48.931 71.007 ;
      RECT 46.401 70.911 48.977 70.961 ;
      RECT 46.447 70.865 49.023 70.915 ;
      RECT 46.493 70.819 49.069 70.869 ;
      RECT 46.539 70.773 49.115 70.823 ;
      RECT 46.585 70.727 49.161 70.777 ;
      RECT 46.631 70.681 49.207 70.731 ;
      RECT 46.677 70.635 49.253 70.685 ;
      RECT 46.723 70.589 49.299 70.639 ;
      RECT 46.769 70.543 49.345 70.593 ;
      RECT 46.815 70.497 49.391 70.547 ;
      RECT 46.861 70.451 49.437 70.501 ;
      RECT 46.907 70.405 49.483 70.455 ;
      RECT 46.953 70.359 49.529 70.409 ;
      RECT 46.999 70.313 49.575 70.363 ;
      RECT 47.045 70.267 49.621 70.317 ;
      RECT 47.091 70.221 49.667 70.271 ;
      RECT 47.137 70.175 49.713 70.225 ;
      RECT 47.183 70.129 49.759 70.179 ;
      RECT 47.229 70.083 49.805 70.133 ;
      RECT 47.275 70.037 49.851 70.087 ;
      RECT 47.321 69.991 49.897 70.041 ;
      RECT 47.367 69.945 49.943 69.995 ;
      RECT 47.413 69.899 49.989 69.949 ;
      RECT 47.459 69.853 50.035 69.903 ;
      RECT 47.505 69.807 50.081 69.857 ;
      RECT 47.551 69.761 50.127 69.811 ;
      RECT 47.597 69.715 50.173 69.765 ;
      RECT 47.643 69.669 50.219 69.719 ;
      RECT 47.689 69.623 50.265 69.673 ;
      RECT 47.735 69.577 50.311 69.627 ;
      RECT 47.781 69.531 50.357 69.581 ;
      RECT 47.827 69.485 50.403 69.535 ;
      RECT 47.873 69.439 50.449 69.489 ;
      RECT 47.919 69.393 50.495 69.443 ;
      RECT 47.965 69.347 50.541 69.397 ;
      RECT 48.011 69.301 50.587 69.351 ;
      RECT 48.057 69.255 50.633 69.305 ;
      RECT 48.103 69.209 50.679 69.259 ;
      RECT 48.149 69.163 50.725 69.213 ;
      RECT 48.195 69.117 50.771 69.167 ;
      RECT 48.241 69.071 50.817 69.121 ;
      RECT 48.287 69.025 50.863 69.075 ;
      RECT 48.333 68.979 50.909 69.029 ;
      RECT 48.379 68.933 50.955 68.983 ;
      RECT 48.425 68.887 51.001 68.937 ;
      RECT 48.471 68.841 51.047 68.891 ;
      RECT 48.517 68.795 51.093 68.845 ;
      RECT 48.563 68.749 51.139 68.799 ;
      RECT 48.609 68.703 51.185 68.753 ;
      RECT 48.655 68.657 51.231 68.707 ;
      RECT 48.701 68.611 51.277 68.661 ;
      RECT 48.747 68.565 51.323 68.615 ;
      RECT 48.793 68.519 51.369 68.569 ;
      RECT 48.839 68.473 51.415 68.523 ;
      RECT 48.885 68.427 51.461 68.477 ;
      RECT 48.931 68.381 51.507 68.431 ;
      RECT 48.977 68.335 51.553 68.385 ;
      RECT 49.023 68.289 51.599 68.339 ;
      RECT 49.069 68.243 51.645 68.293 ;
      RECT 49.115 68.197 51.691 68.247 ;
      RECT 49.161 68.151 51.737 68.201 ;
      RECT 49.207 68.105 51.783 68.155 ;
      RECT 49.253 68.059 51.829 68.109 ;
      RECT 49.299 68.013 51.875 68.063 ;
      RECT 49.345 67.967 51.921 68.017 ;
      RECT 49.391 67.921 51.967 67.971 ;
      RECT 49.437 67.875 52.013 67.925 ;
      RECT 49.483 67.829 52.059 67.879 ;
      RECT 49.529 67.783 52.105 67.833 ;
      RECT 49.575 67.737 52.151 67.787 ;
      RECT 49.621 67.691 52.197 67.741 ;
      RECT 49.667 67.645 52.243 67.695 ;
      RECT 49.713 67.599 52.289 67.649 ;
      RECT 49.759 67.553 52.335 67.603 ;
      RECT 49.805 67.507 52.381 67.557 ;
      RECT 49.851 67.461 52.427 67.511 ;
      RECT 49.897 67.415 52.473 67.465 ;
      RECT 49.943 67.369 52.519 67.419 ;
      RECT 49.989 67.323 52.565 67.373 ;
      RECT 50.035 67.277 52.611 67.327 ;
      RECT 50.081 67.231 52.657 67.281 ;
      RECT 50.127 67.185 52.703 67.235 ;
      RECT 50.173 67.139 52.749 67.189 ;
      RECT 50.219 67.093 52.795 67.143 ;
      RECT 50.265 67.047 52.841 67.097 ;
      RECT 50.311 67.001 52.887 67.051 ;
      RECT 50.357 66.955 52.933 67.005 ;
      RECT 50.403 66.909 52.979 66.959 ;
      RECT 50.449 66.863 53.025 66.913 ;
      RECT 50.495 66.817 53.071 66.867 ;
      RECT 50.541 66.771 53.117 66.821 ;
      RECT 50.587 66.725 53.163 66.775 ;
      RECT 50.633 66.679 53.209 66.729 ;
      RECT 50.679 66.633 53.255 66.683 ;
      RECT 50.725 66.587 53.301 66.637 ;
      RECT 50.771 66.541 53.347 66.591 ;
      RECT 50.817 66.495 53.393 66.545 ;
      RECT 50.863 66.449 53.439 66.499 ;
      RECT 50.909 66.403 53.485 66.453 ;
      RECT 50.955 66.357 53.531 66.407 ;
      RECT 51.001 66.311 53.577 66.361 ;
      RECT 51.047 66.265 53.623 66.315 ;
      RECT 51.093 66.219 53.669 66.269 ;
      RECT 51.139 66.173 53.715 66.223 ;
      RECT 51.185 66.127 53.761 66.177 ;
      RECT 51.231 66.081 53.807 66.131 ;
      RECT 51.277 66.035 53.853 66.085 ;
      RECT 51.323 65.989 53.899 66.039 ;
      RECT 51.369 65.943 53.945 65.993 ;
      RECT 51.415 65.897 53.991 65.947 ;
      RECT 51.461 65.851 54.037 65.901 ;
      RECT 51.507 65.805 54.083 65.855 ;
      RECT 51.553 65.759 54.129 65.809 ;
      RECT 51.599 65.713 54.175 65.763 ;
      RECT 51.645 65.667 54.221 65.717 ;
      RECT 51.691 65.621 54.267 65.671 ;
      RECT 51.737 65.575 54.313 65.625 ;
      RECT 51.783 65.529 54.359 65.579 ;
      RECT 51.829 65.483 54.405 65.533 ;
      RECT 51.875 65.437 54.451 65.487 ;
      RECT 51.921 65.391 54.497 65.441 ;
      RECT 51.967 65.345 54.543 65.395 ;
      RECT 52.013 65.299 54.589 65.349 ;
      RECT 52.059 65.253 54.635 65.303 ;
      RECT 52.105 65.207 54.681 65.257 ;
      RECT 52.151 65.161 54.727 65.211 ;
      RECT 52.197 65.115 54.773 65.165 ;
      RECT 52.243 65.069 54.819 65.119 ;
      RECT 52.289 65.023 54.865 65.073 ;
      RECT 52.335 64.977 54.911 65.027 ;
      RECT 52.381 64.931 54.957 64.981 ;
      RECT 52.427 64.885 55.003 64.935 ;
      RECT 52.473 64.839 55.049 64.889 ;
      RECT 52.519 64.793 55.095 64.843 ;
      RECT 52.565 64.747 55.141 64.797 ;
      RECT 52.611 64.701 55.187 64.751 ;
      RECT 52.657 64.655 55.233 64.705 ;
      RECT 52.703 64.609 55.279 64.659 ;
      RECT 52.749 64.563 55.325 64.613 ;
      RECT 52.795 64.517 55.371 64.567 ;
      RECT 52.841 64.471 55.417 64.521 ;
      RECT 52.887 64.425 55.463 64.475 ;
      RECT 52.933 64.379 55.509 64.429 ;
      RECT 52.979 64.333 55.555 64.383 ;
      RECT 53.025 64.287 55.601 64.337 ;
      RECT 53.071 64.241 55.647 64.291 ;
      RECT 53.117 64.195 55.693 64.245 ;
      RECT 53.163 64.149 55.739 64.199 ;
      RECT 53.209 64.103 55.785 64.153 ;
      RECT 53.255 64.057 55.825 64.11 ;
      RECT 53.301 64.011 55.871 64.067 ;
      RECT 53.347 63.965 55.917 64.021 ;
      RECT 53.393 63.919 55.963 63.975 ;
      RECT 53.439 63.873 56.009 63.929 ;
      RECT 53.485 63.827 56.055 63.883 ;
      RECT 53.531 63.781 56.101 63.837 ;
      RECT 53.577 63.735 56.147 63.791 ;
      RECT 53.623 63.689 56.193 63.745 ;
      RECT 53.669 63.643 56.239 63.699 ;
      RECT 53.715 63.597 56.285 63.653 ;
      RECT 53.761 63.551 56.331 63.607 ;
      RECT 53.807 63.505 56.377 63.561 ;
      RECT 53.853 63.459 56.423 63.515 ;
      RECT 53.899 63.413 56.469 63.469 ;
      RECT 53.945 63.367 56.515 63.423 ;
      RECT 53.991 63.321 56.561 63.377 ;
      RECT 54.037 63.275 56.607 63.331 ;
      RECT 54.083 63.229 56.653 63.285 ;
      RECT 54.129 63.183 56.699 63.239 ;
      RECT 54.175 63.137 56.745 63.193 ;
      RECT 54.221 63.091 56.791 63.147 ;
      RECT 54.267 63.045 56.837 63.101 ;
      RECT 54.313 62.999 56.883 63.055 ;
      RECT 54.359 62.953 56.929 63.009 ;
      RECT 54.405 62.907 56.975 62.963 ;
      RECT 54.451 62.861 57.021 62.917 ;
      RECT 54.497 62.815 57.067 62.871 ;
      RECT 54.543 62.769 57.113 62.825 ;
      RECT 54.589 62.723 57.159 62.779 ;
      RECT 54.635 62.677 57.205 62.733 ;
      RECT 54.681 62.631 57.251 62.687 ;
      RECT 54.727 62.585 57.297 62.641 ;
      RECT 54.773 62.539 57.343 62.595 ;
      RECT 54.819 62.493 57.389 62.549 ;
      RECT 54.865 62.447 57.435 62.503 ;
      RECT 54.911 62.401 57.481 62.457 ;
      RECT 54.957 62.355 57.527 62.411 ;
      RECT 55.003 62.309 57.573 62.365 ;
      RECT 55.049 62.263 57.619 62.319 ;
      RECT 55.095 62.217 57.665 62.273 ;
      RECT 55.141 62.171 57.711 62.227 ;
      RECT 55.187 62.125 57.757 62.181 ;
      RECT 55.233 62.079 57.803 62.135 ;
      RECT 55.279 62.033 57.849 62.089 ;
      RECT 55.325 61.987 57.895 62.043 ;
      RECT 55.371 61.941 57.941 61.997 ;
      RECT 55.417 61.895 57.987 61.951 ;
      RECT 55.463 61.849 58.033 61.905 ;
      RECT 55.509 61.803 58.079 61.859 ;
      RECT 55.555 61.757 58.125 61.813 ;
      RECT 55.601 61.711 58.171 61.767 ;
      RECT 55.647 61.665 58.217 61.721 ;
      RECT 55.693 61.619 58.263 61.675 ;
      RECT 55.739 61.573 58.309 61.629 ;
      RECT 55.785 61.527 58.355 61.583 ;
      RECT 55.831 61.481 58.401 61.537 ;
      RECT 55.877 61.435 58.447 61.491 ;
      RECT 55.923 61.389 58.493 61.445 ;
      RECT 55.969 61.343 58.539 61.399 ;
      RECT 56.015 61.297 58.585 61.353 ;
      RECT 56.061 61.251 58.631 61.307 ;
      RECT 56.107 61.205 58.677 61.261 ;
      RECT 56.153 61.159 58.723 61.215 ;
      RECT 56.199 61.113 58.769 61.169 ;
      RECT 56.245 61.067 58.815 61.123 ;
      RECT 56.291 61.021 58.861 61.077 ;
      RECT 56.337 60.975 58.907 61.031 ;
      RECT 56.383 60.929 58.953 60.985 ;
      RECT 56.429 60.883 58.999 60.939 ;
      RECT 56.475 60.837 59.045 60.893 ;
      RECT 56.521 60.791 59.091 60.847 ;
      RECT 56.567 60.745 59.137 60.801 ;
      RECT 56.613 60.699 59.183 60.755 ;
      RECT 56.659 60.653 59.229 60.709 ;
      RECT 56.705 60.607 59.275 60.663 ;
      RECT 56.751 60.561 59.321 60.617 ;
      RECT 56.797 60.515 59.367 60.571 ;
      RECT 56.843 60.469 59.413 60.525 ;
      RECT 56.889 60.423 59.459 60.479 ;
      RECT 56.935 60.377 59.505 60.433 ;
      RECT 56.981 60.331 59.551 60.387 ;
      RECT 57.027 60.285 59.597 60.341 ;
      RECT 57.073 60.239 59.643 60.295 ;
      RECT 57.119 60.193 59.689 60.249 ;
      RECT 57.165 60.147 59.735 60.203 ;
      RECT 57.211 60.101 59.781 60.157 ;
      RECT 57.257 60.055 59.827 60.111 ;
      RECT 57.303 60.009 59.873 60.065 ;
      RECT 57.349 59.963 59.919 60.019 ;
      RECT 57.395 59.917 59.965 59.973 ;
      RECT 57.441 59.871 60.011 59.927 ;
      RECT 57.487 59.825 60.057 59.881 ;
      RECT 57.533 59.779 60.103 59.835 ;
      RECT 57.579 59.733 60.149 59.789 ;
      RECT 57.625 59.687 60.195 59.743 ;
      RECT 57.671 59.641 60.241 59.697 ;
      RECT 57.717 59.595 60.287 59.651 ;
      RECT 57.763 59.549 60.333 59.605 ;
      RECT 57.809 59.503 60.379 59.559 ;
      RECT 57.855 59.457 60.425 59.513 ;
      RECT 57.901 59.411 60.471 59.467 ;
      RECT 57.947 59.365 60.517 59.421 ;
      RECT 57.993 59.319 60.563 59.375 ;
      RECT 58.039 59.273 60.609 59.329 ;
      RECT 58.085 59.227 60.655 59.283 ;
      RECT 58.131 59.181 60.701 59.237 ;
      RECT 58.177 59.135 60.747 59.191 ;
      RECT 58.223 59.089 60.793 59.145 ;
      RECT 58.269 59.043 60.839 59.099 ;
      RECT 58.315 58.997 60.885 59.053 ;
      RECT 58.361 58.951 60.931 59.007 ;
      RECT 58.407 58.905 60.977 58.961 ;
      RECT 58.453 58.859 61.023 58.915 ;
      RECT 58.499 58.813 61.069 58.869 ;
      RECT 58.545 58.767 61.115 58.823 ;
      RECT 58.591 58.721 61.161 58.777 ;
      RECT 58.637 58.675 61.207 58.731 ;
      RECT 58.683 58.629 61.253 58.685 ;
      RECT 58.729 58.583 61.299 58.639 ;
      RECT 58.775 58.537 61.345 58.593 ;
      RECT 58.821 58.491 61.391 58.547 ;
      RECT 58.867 58.445 61.437 58.501 ;
      RECT 58.913 58.399 61.483 58.455 ;
      RECT 58.959 58.353 61.529 58.409 ;
      RECT 59.005 58.307 61.575 58.363 ;
      RECT 59.051 58.261 61.621 58.317 ;
      RECT 59.097 58.215 61.667 58.271 ;
      RECT 59.143 58.169 61.713 58.225 ;
      RECT 59.189 58.123 61.759 58.179 ;
      RECT 59.235 58.077 61.805 58.133 ;
      RECT 59.281 58.031 61.851 58.087 ;
      RECT 59.327 57.985 61.897 58.041 ;
      RECT 59.373 57.939 61.943 57.995 ;
      RECT 59.419 57.893 61.989 57.949 ;
      RECT 59.465 57.847 62.035 57.903 ;
      RECT 59.511 57.801 62.081 57.857 ;
      RECT 59.557 57.755 62.127 57.811 ;
      RECT 59.603 57.709 62.173 57.765 ;
      RECT 59.649 57.663 62.219 57.719 ;
      RECT 59.695 57.617 62.265 57.673 ;
      RECT 59.741 57.571 62.311 57.627 ;
      RECT 59.787 57.525 62.357 57.581 ;
      RECT 59.833 57.479 62.403 57.535 ;
      RECT 59.879 57.433 62.449 57.489 ;
      RECT 59.925 57.387 62.495 57.443 ;
      RECT 59.971 57.341 62.541 57.397 ;
      RECT 60.017 57.295 62.587 57.351 ;
      RECT 60.063 57.249 62.633 57.305 ;
      RECT 60.109 57.203 62.679 57.259 ;
      RECT 60.155 57.157 62.725 57.213 ;
      RECT 60.201 57.111 62.771 57.167 ;
      RECT 60.247 57.065 62.817 57.121 ;
      RECT 60.293 57.019 62.863 57.075 ;
      RECT 60.339 56.973 62.909 57.029 ;
      RECT 60.385 56.927 62.955 56.983 ;
      RECT 60.431 56.881 63.001 56.937 ;
      RECT 60.477 56.835 63.047 56.891 ;
      RECT 60.523 56.789 63.093 56.845 ;
      RECT 60.569 56.743 63.139 56.799 ;
      RECT 60.615 56.697 63.185 56.753 ;
      RECT 60.661 56.651 63.231 56.707 ;
      RECT 60.707 56.605 63.277 56.661 ;
      RECT 60.753 56.559 63.323 56.615 ;
      RECT 60.799 56.513 63.369 56.569 ;
      RECT 60.845 56.467 63.415 56.523 ;
      RECT 60.891 56.421 63.461 56.477 ;
      RECT 60.937 56.375 63.507 56.431 ;
      RECT 60.983 56.329 63.553 56.385 ;
      RECT 61.029 56.283 63.599 56.339 ;
      RECT 61.075 56.237 63.645 56.293 ;
      RECT 61.121 56.191 63.691 56.247 ;
      RECT 61.167 56.145 63.737 56.201 ;
      RECT 61.213 56.099 63.783 56.155 ;
      RECT 61.259 56.053 63.829 56.109 ;
      RECT 61.305 56.007 63.875 56.063 ;
      RECT 61.351 55.961 63.921 56.017 ;
      RECT 61.397 55.915 63.967 55.971 ;
      RECT 61.443 55.869 64.013 55.925 ;
      RECT 61.489 55.823 64.059 55.879 ;
      RECT 61.535 55.777 64.105 55.833 ;
      RECT 61.581 55.731 64.151 55.787 ;
      RECT 61.627 55.685 64.197 55.741 ;
      RECT 61.673 55.639 64.243 55.695 ;
      RECT 61.719 55.593 64.289 55.649 ;
      RECT 61.765 55.547 64.335 55.603 ;
      RECT 61.811 55.501 64.381 55.557 ;
      RECT 61.857 55.455 64.427 55.511 ;
      RECT 61.903 55.409 64.473 55.465 ;
      RECT 61.949 55.363 64.519 55.419 ;
      RECT 61.995 55.317 64.565 55.373 ;
      RECT 62.041 55.271 64.611 55.327 ;
      RECT 62.087 55.225 64.657 55.281 ;
      RECT 62.133 55.179 64.703 55.235 ;
      RECT 62.179 55.133 64.749 55.189 ;
      RECT 62.225 55.087 64.795 55.143 ;
      RECT 62.271 55.041 64.841 55.097 ;
      RECT 62.317 54.995 64.887 55.051 ;
      RECT 62.363 54.949 64.933 55.005 ;
      RECT 62.409 54.903 64.979 54.959 ;
      RECT 62.455 54.857 65.025 54.913 ;
      RECT 62.501 54.811 65.071 54.867 ;
      RECT 62.547 54.765 65.117 54.821 ;
      RECT 62.593 54.719 65.163 54.775 ;
      RECT 62.639 54.673 65.209 54.729 ;
      RECT 62.685 54.627 65.255 54.683 ;
      RECT 62.731 54.581 65.301 54.637 ;
      RECT 62.777 54.535 65.347 54.591 ;
      RECT 62.823 54.489 65.393 54.545 ;
      RECT 62.869 54.443 65.439 54.499 ;
      RECT 62.915 54.397 65.485 54.453 ;
      RECT 62.961 54.351 65.531 54.407 ;
      RECT 63.007 54.305 65.577 54.361 ;
      RECT 63.053 54.259 65.623 54.315 ;
      RECT 63.099 54.213 65.669 54.269 ;
      RECT 63.145 54.167 65.715 54.223 ;
      RECT 63.191 54.121 65.761 54.177 ;
      RECT 63.237 54.075 65.807 54.131 ;
      RECT 63.283 54.029 65.853 54.085 ;
      RECT 63.329 53.983 65.899 54.039 ;
      RECT 63.375 53.937 65.945 53.993 ;
      RECT 63.421 53.891 65.991 53.947 ;
      RECT 63.467 53.845 66.037 53.901 ;
      RECT 63.513 53.799 66.083 53.855 ;
      RECT 63.559 53.753 66.129 53.809 ;
      RECT 63.605 53.707 66.175 53.763 ;
      RECT 63.651 53.661 66.221 53.717 ;
      RECT 63.697 53.615 66.267 53.671 ;
      RECT 63.743 53.569 66.313 53.625 ;
      RECT 63.789 53.523 66.359 53.579 ;
      RECT 63.835 53.477 66.405 53.533 ;
      RECT 63.881 53.431 66.451 53.487 ;
      RECT 63.927 53.385 66.497 53.441 ;
      RECT 63.973 53.339 66.543 53.395 ;
      RECT 64.019 53.293 66.589 53.349 ;
      RECT 64.065 53.247 66.635 53.303 ;
      RECT 64.111 53.201 66.681 53.257 ;
      RECT 64.157 53.155 66.727 53.211 ;
      RECT 64.203 53.109 66.773 53.165 ;
      RECT 64.249 53.063 66.819 53.119 ;
      RECT 64.295 53.017 66.865 53.073 ;
      RECT 64.341 52.971 66.911 53.027 ;
      RECT 64.387 52.925 66.957 52.981 ;
      RECT 64.433 52.879 67.003 52.935 ;
      RECT 64.479 52.833 67.049 52.889 ;
      RECT 64.525 52.787 67.095 52.843 ;
      RECT 64.571 52.741 67.141 52.797 ;
      RECT 64.617 52.695 67.187 52.751 ;
      RECT 64.663 52.649 67.233 52.705 ;
      RECT 64.709 52.603 67.279 52.659 ;
      RECT 64.755 52.557 67.325 52.613 ;
      RECT 64.801 52.511 67.371 52.567 ;
      RECT 64.847 52.465 67.417 52.521 ;
      RECT 64.893 52.419 67.463 52.475 ;
      RECT 64.939 52.373 67.509 52.429 ;
      RECT 64.985 52.327 67.555 52.383 ;
      RECT 65.031 52.281 67.601 52.337 ;
      RECT 65.077 52.235 67.647 52.291 ;
      RECT 65.123 52.189 67.693 52.245 ;
      RECT 65.169 52.143 67.739 52.199 ;
      RECT 65.215 52.097 67.785 52.153 ;
      RECT 65.261 52.051 67.831 52.107 ;
      RECT 65.307 52.005 67.877 52.061 ;
      RECT 65.353 51.959 67.923 52.015 ;
      RECT 65.399 51.913 67.969 51.969 ;
      RECT 65.445 51.867 68.015 51.923 ;
      RECT 65.491 51.821 68.061 51.877 ;
      RECT 65.537 51.775 68.107 51.831 ;
      RECT 65.583 51.729 68.153 51.785 ;
      RECT 65.629 51.683 68.199 51.739 ;
      RECT 65.675 51.637 68.245 51.693 ;
      RECT 65.721 51.591 68.291 51.647 ;
      RECT 65.767 51.545 68.337 51.601 ;
      RECT 65.813 51.499 68.383 51.555 ;
      RECT 65.859 51.453 68.429 51.509 ;
      RECT 65.905 51.407 68.475 51.463 ;
      RECT 65.951 51.361 68.521 51.417 ;
      RECT 65.997 51.315 68.567 51.371 ;
      RECT 66.043 51.269 68.613 51.325 ;
      RECT 66.089 51.223 68.659 51.279 ;
      RECT 66.135 51.177 68.705 51.233 ;
      RECT 66.181 51.131 68.751 51.187 ;
      RECT 66.227 51.085 68.797 51.141 ;
      RECT 66.273 51.039 68.843 51.095 ;
      RECT 66.319 50.993 68.889 51.049 ;
      RECT 66.365 50.947 68.935 51.003 ;
      RECT 66.411 50.901 68.981 50.957 ;
      RECT 66.457 50.855 69.027 50.911 ;
      RECT 66.503 50.809 69.073 50.865 ;
      RECT 66.549 50.763 69.119 50.819 ;
      RECT 66.595 50.717 69.165 50.773 ;
      RECT 66.641 50.671 69.211 50.727 ;
      RECT 66.687 50.625 69.257 50.681 ;
      RECT 66.733 50.579 69.303 50.635 ;
      RECT 66.779 50.533 69.349 50.589 ;
      RECT 66.825 50.487 69.395 50.543 ;
      RECT 66.871 50.441 69.441 50.497 ;
      RECT 66.917 50.395 69.487 50.451 ;
      RECT 66.963 50.349 69.533 50.405 ;
      RECT 67.009 50.303 69.579 50.359 ;
      RECT 67.055 50.257 69.625 50.313 ;
      RECT 67.101 50.211 69.671 50.267 ;
      RECT 67.147 50.165 69.717 50.221 ;
      RECT 69.677 47.652 69.717 50.221 ;
      RECT 67.193 50.119 69.763 50.175 ;
      RECT 69.69 47.622 69.763 50.175 ;
      RECT 67.239 50.073 69.809 50.129 ;
      RECT 69.736 47.576 69.809 50.129 ;
      RECT 67.285 50.027 69.855 50.083 ;
      RECT 69.782 47.53 69.855 50.083 ;
      RECT 67.331 49.981 69.901 50.037 ;
      RECT 69.828 47.484 69.901 50.037 ;
      RECT 67.377 49.935 69.947 49.991 ;
      RECT 69.874 47.438 69.947 49.991 ;
      RECT 67.423 49.889 69.993 49.945 ;
      RECT 69.92 47.392 69.993 49.945 ;
      RECT 67.469 49.843 70.039 49.899 ;
      RECT 69.966 47.346 70.039 49.899 ;
      RECT 67.515 49.797 70.085 49.853 ;
      RECT 70.012 47.3 70.085 49.853 ;
      RECT 67.561 49.751 70.131 49.807 ;
      RECT 70.058 47.254 70.131 49.807 ;
      RECT 67.607 49.705 70.177 49.761 ;
      RECT 70.104 47.208 70.177 49.761 ;
      RECT 67.653 49.659 70.223 49.715 ;
      RECT 70.15 47.162 70.223 49.715 ;
      RECT 67.699 49.613 70.269 49.669 ;
      RECT 70.196 47.116 70.269 49.669 ;
      RECT 67.745 49.567 70.315 49.623 ;
      RECT 70.242 47.07 70.315 49.623 ;
      RECT 67.791 49.521 70.361 49.577 ;
      RECT 70.288 47.024 70.361 49.577 ;
      RECT 67.837 49.475 70.407 49.531 ;
      RECT 70.334 46.978 70.407 49.531 ;
      RECT 67.883 49.429 70.453 49.485 ;
      RECT 70.38 46.932 70.453 49.485 ;
      RECT 67.929 49.383 70.499 49.439 ;
      RECT 70.426 46.886 70.499 49.439 ;
      RECT 67.975 49.337 70.545 49.393 ;
      RECT 70.472 46.84 70.545 49.393 ;
      RECT 68.021 49.291 70.591 49.347 ;
      RECT 70.518 46.794 70.591 49.347 ;
      RECT 68.067 49.245 70.637 49.301 ;
      RECT 70.564 46.748 70.637 49.301 ;
      RECT 68.113 49.199 70.683 49.255 ;
      RECT 70.61 46.702 70.683 49.255 ;
      RECT 68.159 49.153 70.729 49.209 ;
      RECT 70.656 46.656 70.729 49.209 ;
      RECT 68.205 49.107 70.775 49.163 ;
      RECT 70.702 46.61 70.775 49.163 ;
      RECT 68.251 49.061 70.821 49.117 ;
      RECT 70.748 46.564 70.821 49.117 ;
      RECT 68.297 49.015 70.867 49.071 ;
      RECT 70.794 46.518 70.867 49.071 ;
      RECT 68.343 48.969 70.913 49.025 ;
      RECT 70.84 46.472 70.913 49.025 ;
      RECT 68.389 48.923 70.959 48.979 ;
      RECT 70.886 46.426 70.959 48.979 ;
      RECT 68.435 48.877 71.005 48.933 ;
      RECT 70.932 46.38 71.005 48.933 ;
      RECT 68.481 48.831 71.051 48.887 ;
      RECT 70.978 46.334 71.051 48.887 ;
      RECT 68.527 48.785 71.097 48.841 ;
      RECT 71.024 46.288 71.097 48.841 ;
      RECT 68.573 48.739 71.143 48.795 ;
      RECT 71.07 46.242 71.143 48.795 ;
      RECT 68.619 48.693 71.189 48.749 ;
      RECT 71.116 46.196 71.189 48.749 ;
      RECT 68.665 48.647 71.235 48.703 ;
      RECT 71.162 46.15 71.235 48.703 ;
      RECT 68.711 48.601 71.281 48.657 ;
      RECT 71.208 46.104 71.281 48.657 ;
      RECT 68.757 48.555 71.327 48.611 ;
      RECT 71.254 46.058 71.327 48.611 ;
      RECT 68.803 48.509 71.373 48.565 ;
      RECT 71.3 46.012 71.373 48.565 ;
      RECT 68.849 48.463 71.419 48.519 ;
      RECT 71.346 45.966 71.419 48.519 ;
      RECT 68.895 48.417 71.465 48.473 ;
      RECT 71.392 45.92 71.465 48.473 ;
      RECT 68.941 48.371 71.511 48.427 ;
      RECT 71.438 45.874 71.511 48.427 ;
      RECT 68.987 48.325 71.557 48.381 ;
      RECT 71.484 45.828 71.557 48.381 ;
      RECT 69.033 48.279 71.603 48.335 ;
      RECT 71.53 45.782 71.603 48.335 ;
      RECT 69.079 48.233 71.649 48.289 ;
      RECT 71.576 45.736 71.649 48.289 ;
      RECT 69.125 48.187 71.695 48.243 ;
      RECT 71.622 45.69 71.695 48.243 ;
      RECT 69.171 48.141 71.741 48.197 ;
      RECT 71.668 45.644 71.741 48.197 ;
      RECT 69.217 48.095 71.787 48.151 ;
      RECT 71.714 45.598 71.787 48.151 ;
      RECT 69.263 48.049 71.833 48.105 ;
      RECT 71.76 45.552 71.833 48.105 ;
      RECT 69.309 48.003 71.879 48.059 ;
      RECT 71.806 45.506 71.879 48.059 ;
      RECT 69.355 47.957 71.925 48.013 ;
      RECT 71.852 45.46 71.925 48.013 ;
      RECT 69.401 47.911 71.971 47.967 ;
      RECT 71.898 45.414 71.971 47.967 ;
      RECT 69.447 47.865 72.017 47.921 ;
      RECT 71.944 45.368 72.017 47.921 ;
      RECT 69.493 47.819 72.063 47.875 ;
      RECT 71.99 45.322 72.063 47.875 ;
      RECT 69.539 47.773 72.109 47.829 ;
      RECT 72.036 45.276 72.109 47.829 ;
      RECT 69.585 47.727 72.155 47.783 ;
      RECT 72.082 45.23 72.155 47.783 ;
      RECT 69.631 47.681 72.201 47.737 ;
      RECT 72.128 45.184 72.201 47.737 ;
      RECT 72.174 45.138 72.247 47.691 ;
      RECT 72.22 45.092 72.293 47.645 ;
      RECT 72.266 45.046 72.339 47.599 ;
      RECT 72.312 45 72.385 47.553 ;
      RECT 72.358 44.954 72.431 47.507 ;
      RECT 72.404 44.908 72.477 47.461 ;
      RECT 72.45 44.862 72.523 47.415 ;
      RECT 72.496 44.816 72.569 47.369 ;
      RECT 72.542 44.77 72.615 47.323 ;
      RECT 72.588 44.724 72.661 47.277 ;
      RECT 72.634 44.678 72.707 47.231 ;
      RECT 72.68 44.632 72.753 47.185 ;
      RECT 72.726 44.586 72.799 47.139 ;
      RECT 72.772 44.54 72.845 47.093 ;
      RECT 72.818 44.494 72.891 47.047 ;
      RECT 72.864 44.448 72.937 47.001 ;
      RECT 72.91 44.402 72.983 46.955 ;
      RECT 72.956 44.356 73.029 46.909 ;
      RECT 73.002 44.31 73.075 46.863 ;
      RECT 73.048 44.264 73.121 46.817 ;
      RECT 73.094 44.218 73.167 46.771 ;
      RECT 73.14 44.172 73.213 46.725 ;
      RECT 73.186 44.126 73.259 46.679 ;
      RECT 73.232 44.08 73.305 46.633 ;
      RECT 73.278 44.034 73.351 46.587 ;
      RECT 73.324 43.988 73.397 46.541 ;
      RECT 73.37 43.942 73.443 46.495 ;
      RECT 73.416 43.896 73.489 46.449 ;
      RECT 73.462 43.85 73.535 46.403 ;
      RECT 73.508 43.804 73.581 46.357 ;
      RECT 73.554 43.758 73.627 46.311 ;
      RECT 73.6 43.712 73.673 46.265 ;
      RECT 73.646 43.666 73.719 46.219 ;
      RECT 73.692 43.62 73.765 46.173 ;
      RECT 73.738 43.574 73.811 46.127 ;
      RECT 73.784 43.528 73.857 46.081 ;
      RECT 73.83 43.482 73.903 46.035 ;
      RECT 73.876 43.436 73.949 45.989 ;
      RECT 73.922 43.39 73.995 45.943 ;
      RECT 73.968 43.344 74.041 45.897 ;
      RECT 74.014 43.298 74.087 45.851 ;
      RECT 74.06 43.252 74.133 45.805 ;
      RECT 74.106 43.206 74.179 45.759 ;
      RECT 74.152 43.16 74.225 45.713 ;
      RECT 74.198 43.114 74.271 45.667 ;
      RECT 74.244 43.068 74.317 45.621 ;
      RECT 74.29 43.022 74.363 45.575 ;
      RECT 74.336 42.976 74.409 45.529 ;
      RECT 74.382 42.93 74.455 45.483 ;
      RECT 74.428 42.884 74.501 45.437 ;
      RECT 74.474 42.838 74.547 45.391 ;
      RECT 74.52 42.792 74.593 45.345 ;
      RECT 74.566 42.746 74.639 45.299 ;
      RECT 74.612 42.699 74.685 45.253 ;
      RECT 74.658 42.675 74.731 45.207 ;
      RECT 74.658 42.675 74.777 45.161 ;
      RECT 74.658 42.675 74.823 45.115 ;
      RECT 74.658 42.675 74.869 45.069 ;
      RECT 74.658 42.675 74.915 45.023 ;
      RECT 74.658 42.675 74.961 44.977 ;
      RECT 74.658 42.675 75.007 44.931 ;
      RECT 74.658 42.675 75.053 44.885 ;
      RECT 74.658 42.675 75.099 44.839 ;
      RECT 74.658 42.675 75.145 44.793 ;
      RECT 74.658 42.675 75.191 44.747 ;
      RECT 74.658 42.675 75.237 44.701 ;
      RECT 74.658 42.675 75.283 44.655 ;
      RECT 74.658 42.675 75.329 44.609 ;
      RECT 74.658 42.675 75.375 44.563 ;
      RECT 74.658 42.675 75.421 44.517 ;
      RECT 74.658 42.675 75.467 44.471 ;
      RECT 74.658 42.675 75.513 44.425 ;
      RECT 74.658 42.675 75.559 44.379 ;
      RECT 74.658 42.675 75.605 44.333 ;
      RECT 74.658 42.675 75.651 44.287 ;
      RECT 74.658 42.675 75.697 44.241 ;
      RECT 74.658 42.675 75.743 44.195 ;
      RECT 74.658 42.675 75.789 44.149 ;
      RECT 74.658 42.675 75.835 44.103 ;
      RECT 74.658 42.675 75.881 44.057 ;
      RECT 74.658 42.675 75.927 44.011 ;
      RECT 74.658 42.675 75.973 43.965 ;
      RECT 74.658 42.675 76.019 43.919 ;
      RECT 74.658 42.675 76.065 43.873 ;
      RECT 73.508 43.804 76.09 43.837 ;
      RECT 74.658 42.675 110 43.825 ;
      RECT 56.175 81.387 57.325 110 ;
      RECT 56.175 81.387 57.371 82.562 ;
      RECT 56.175 81.387 57.417 82.516 ;
      RECT 56.175 81.387 57.463 82.47 ;
      RECT 56.175 81.387 57.509 82.424 ;
      RECT 56.175 81.387 57.555 82.378 ;
      RECT 56.175 81.387 57.601 82.332 ;
      RECT 56.175 81.387 57.647 82.286 ;
      RECT 56.175 81.387 57.693 82.24 ;
      RECT 56.175 81.387 57.739 82.194 ;
      RECT 56.175 81.387 57.785 82.148 ;
      RECT 56.175 81.387 57.831 82.102 ;
      RECT 56.175 81.387 57.877 82.056 ;
      RECT 56.175 81.387 57.923 82.01 ;
      RECT 56.175 81.387 57.969 81.964 ;
      RECT 56.175 81.387 58.015 81.918 ;
      RECT 56.175 81.387 58.061 81.872 ;
      RECT 56.175 81.387 58.107 81.826 ;
      RECT 56.175 81.387 58.153 81.78 ;
      RECT 56.175 81.387 58.199 81.734 ;
      RECT 56.175 81.387 58.245 81.688 ;
      RECT 56.175 81.387 58.291 81.642 ;
      RECT 56.175 81.387 58.337 81.596 ;
      RECT 56.175 81.387 58.383 81.55 ;
      RECT 56.175 81.387 58.429 81.504 ;
      RECT 56.175 81.387 58.475 81.458 ;
      RECT 56.221 81.341 58.521 81.412 ;
      RECT 56.267 81.295 58.567 81.366 ;
      RECT 56.313 81.249 58.613 81.32 ;
      RECT 56.359 81.203 58.659 81.274 ;
      RECT 56.405 81.157 58.705 81.228 ;
      RECT 56.451 81.111 58.751 81.182 ;
      RECT 56.497 81.065 58.797 81.136 ;
      RECT 56.543 81.019 58.843 81.09 ;
      RECT 56.589 80.973 58.889 81.044 ;
      RECT 56.635 80.927 58.935 80.998 ;
      RECT 56.681 80.881 58.981 80.952 ;
      RECT 56.727 80.835 59.027 80.906 ;
      RECT 56.773 80.789 59.073 80.86 ;
      RECT 56.819 80.743 59.119 80.814 ;
      RECT 56.865 80.697 59.165 80.768 ;
      RECT 56.911 80.651 59.211 80.722 ;
      RECT 56.957 80.605 59.257 80.676 ;
      RECT 57.003 80.559 59.303 80.63 ;
      RECT 57.049 80.513 59.349 80.584 ;
      RECT 57.095 80.467 59.395 80.538 ;
      RECT 57.141 80.421 59.441 80.492 ;
      RECT 57.187 80.375 59.487 80.446 ;
      RECT 57.233 80.329 59.533 80.4 ;
      RECT 57.279 80.283 59.579 80.354 ;
      RECT 57.325 80.237 59.625 80.308 ;
      RECT 57.371 80.191 59.671 80.262 ;
      RECT 57.417 80.145 59.717 80.216 ;
      RECT 57.463 80.099 59.763 80.17 ;
      RECT 57.509 80.053 59.809 80.124 ;
      RECT 57.555 80.007 59.855 80.078 ;
      RECT 57.601 79.961 59.901 80.032 ;
      RECT 57.647 79.915 59.947 79.986 ;
      RECT 57.693 79.869 59.993 79.94 ;
      RECT 57.739 79.823 60.039 79.894 ;
      RECT 57.785 79.777 60.085 79.848 ;
      RECT 57.831 79.731 60.131 79.802 ;
      RECT 57.877 79.685 60.177 79.756 ;
      RECT 57.923 79.639 60.223 79.71 ;
      RECT 57.969 79.593 60.269 79.664 ;
      RECT 58.015 79.547 60.315 79.618 ;
      RECT 58.061 79.501 60.361 79.572 ;
      RECT 58.107 79.455 60.407 79.526 ;
      RECT 58.153 79.409 60.453 79.48 ;
      RECT 58.199 79.363 60.499 79.434 ;
      RECT 58.245 79.317 60.545 79.388 ;
      RECT 58.291 79.271 60.591 79.342 ;
      RECT 58.337 79.225 60.637 79.296 ;
      RECT 58.383 79.179 60.683 79.25 ;
      RECT 58.429 79.133 60.729 79.204 ;
      RECT 58.475 79.087 60.775 79.158 ;
      RECT 58.521 79.041 60.821 79.112 ;
      RECT 58.567 78.995 60.867 79.066 ;
      RECT 58.613 78.949 60.913 79.02 ;
      RECT 58.659 78.903 60.959 78.974 ;
      RECT 58.705 78.857 61.005 78.928 ;
      RECT 58.751 78.811 61.051 78.882 ;
      RECT 58.797 78.765 61.097 78.836 ;
      RECT 58.843 78.719 61.143 78.79 ;
      RECT 58.889 78.673 61.189 78.744 ;
      RECT 58.935 78.627 61.235 78.698 ;
      RECT 58.981 78.581 61.281 78.652 ;
      RECT 59.027 78.535 61.327 78.606 ;
      RECT 59.073 78.489 61.373 78.56 ;
      RECT 59.119 78.443 61.419 78.514 ;
      RECT 59.165 78.397 61.465 78.468 ;
      RECT 59.211 78.351 61.511 78.422 ;
      RECT 59.257 78.305 61.557 78.376 ;
      RECT 59.303 78.259 61.603 78.33 ;
      RECT 59.349 78.213 61.649 78.284 ;
      RECT 59.395 78.167 61.695 78.238 ;
      RECT 59.441 78.121 61.741 78.192 ;
      RECT 59.487 78.075 61.787 78.146 ;
      RECT 59.533 78.029 61.833 78.1 ;
      RECT 59.579 77.983 61.879 78.054 ;
      RECT 59.625 77.937 61.925 78.008 ;
      RECT 59.671 77.891 61.971 77.962 ;
      RECT 59.717 77.845 62.017 77.916 ;
      RECT 59.763 77.799 62.063 77.87 ;
      RECT 59.809 77.753 62.109 77.824 ;
      RECT 59.855 77.707 62.155 77.778 ;
      RECT 59.901 77.661 62.201 77.732 ;
      RECT 59.947 77.615 62.247 77.686 ;
      RECT 59.993 77.569 62.293 77.64 ;
      RECT 60.039 77.523 62.339 77.594 ;
      RECT 60.085 77.477 62.385 77.548 ;
      RECT 60.131 77.431 62.431 77.502 ;
      RECT 60.177 77.385 62.477 77.456 ;
      RECT 60.223 77.339 62.523 77.41 ;
      RECT 60.269 77.293 62.569 77.364 ;
      RECT 60.315 77.247 62.615 77.318 ;
      RECT 60.361 77.201 62.661 77.272 ;
      RECT 60.407 77.155 62.707 77.226 ;
      RECT 60.453 77.109 62.753 77.18 ;
      RECT 60.499 77.063 62.799 77.134 ;
      RECT 60.545 77.017 62.845 77.088 ;
      RECT 60.591 76.971 62.891 77.042 ;
      RECT 60.637 76.925 62.937 76.996 ;
      RECT 60.683 76.879 62.983 76.95 ;
      RECT 60.729 76.833 63.029 76.904 ;
      RECT 60.775 76.787 63.075 76.858 ;
      RECT 60.821 76.741 63.121 76.812 ;
      RECT 60.867 76.695 63.167 76.766 ;
      RECT 60.913 76.649 63.213 76.72 ;
      RECT 60.959 76.603 63.259 76.674 ;
      RECT 61.005 76.557 63.305 76.628 ;
      RECT 61.005 76.557 63.325 76.595 ;
      RECT 61.051 76.511 63.371 76.562 ;
      RECT 63.305 74.257 63.371 76.562 ;
      RECT 61.097 76.465 63.417 76.516 ;
      RECT 63.351 74.211 63.417 76.516 ;
      RECT 61.143 76.419 63.463 76.47 ;
      RECT 63.397 74.165 63.463 76.47 ;
      RECT 61.189 76.373 63.509 76.424 ;
      RECT 63.443 74.119 63.509 76.424 ;
      RECT 61.235 76.327 63.555 76.378 ;
      RECT 63.489 74.073 63.555 76.378 ;
      RECT 61.281 76.281 63.601 76.332 ;
      RECT 63.535 74.027 63.601 76.332 ;
      RECT 61.327 76.235 63.647 76.286 ;
      RECT 63.581 73.981 63.647 76.286 ;
      RECT 61.373 76.189 63.693 76.24 ;
      RECT 63.627 73.935 63.693 76.24 ;
      RECT 61.419 76.143 63.739 76.194 ;
      RECT 63.673 73.889 63.739 76.194 ;
      RECT 61.465 76.097 63.785 76.148 ;
      RECT 63.719 73.843 63.785 76.148 ;
      RECT 61.511 76.051 63.831 76.102 ;
      RECT 63.765 73.797 63.831 76.102 ;
      RECT 61.557 76.005 63.877 76.056 ;
      RECT 63.811 73.751 63.877 76.056 ;
      RECT 61.603 75.959 63.923 76.01 ;
      RECT 63.857 73.705 63.923 76.01 ;
      RECT 61.649 75.913 63.969 75.964 ;
      RECT 63.903 73.659 63.969 75.964 ;
      RECT 61.695 75.867 64.015 75.918 ;
      RECT 63.949 73.613 64.015 75.918 ;
      RECT 61.741 75.821 64.061 75.872 ;
      RECT 63.995 73.567 64.061 75.872 ;
      RECT 61.787 75.775 64.107 75.826 ;
      RECT 64.041 73.521 64.107 75.826 ;
      RECT 61.833 75.729 64.153 75.78 ;
      RECT 64.087 73.475 64.153 75.78 ;
      RECT 61.879 75.683 64.199 75.734 ;
      RECT 64.133 73.429 64.199 75.734 ;
      RECT 61.925 75.637 64.245 75.688 ;
      RECT 64.179 73.383 64.245 75.688 ;
      RECT 61.971 75.591 64.291 75.642 ;
      RECT 64.225 73.337 64.291 75.642 ;
      RECT 62.017 75.545 64.337 75.596 ;
      RECT 64.271 73.291 64.337 75.596 ;
      RECT 62.063 75.499 64.383 75.55 ;
      RECT 64.317 73.245 64.383 75.55 ;
      RECT 62.109 75.453 64.429 75.504 ;
      RECT 64.363 73.199 64.429 75.504 ;
      RECT 62.155 75.407 64.475 75.458 ;
      RECT 64.409 73.153 64.475 75.458 ;
      RECT 62.201 75.361 64.521 75.412 ;
      RECT 64.455 73.107 64.521 75.412 ;
      RECT 62.247 75.315 64.567 75.366 ;
      RECT 64.501 73.061 64.567 75.366 ;
      RECT 62.293 75.269 64.613 75.32 ;
      RECT 64.547 73.015 64.613 75.32 ;
      RECT 62.339 75.223 64.659 75.274 ;
      RECT 64.593 72.969 64.659 75.274 ;
      RECT 62.385 75.177 64.705 75.228 ;
      RECT 64.639 72.923 64.705 75.228 ;
      RECT 62.431 75.131 64.751 75.182 ;
      RECT 64.685 72.877 64.751 75.182 ;
      RECT 62.477 75.085 64.797 75.136 ;
      RECT 64.731 72.831 64.797 75.136 ;
      RECT 62.523 75.039 64.843 75.09 ;
      RECT 64.777 72.785 64.843 75.09 ;
      RECT 62.569 74.993 64.889 75.044 ;
      RECT 64.823 72.739 64.889 75.044 ;
      RECT 62.615 74.947 64.935 74.998 ;
      RECT 64.869 72.693 64.935 74.998 ;
      RECT 62.661 74.901 64.981 74.952 ;
      RECT 64.915 72.647 64.981 74.952 ;
      RECT 62.707 74.855 65.027 74.906 ;
      RECT 64.961 72.601 65.027 74.906 ;
      RECT 62.753 74.809 65.073 74.86 ;
      RECT 65.007 72.555 65.073 74.86 ;
      RECT 62.799 74.763 65.119 74.814 ;
      RECT 65.053 72.509 65.119 74.814 ;
      RECT 62.845 74.717 65.165 74.768 ;
      RECT 65.099 72.463 65.165 74.768 ;
      RECT 62.891 74.671 65.211 74.722 ;
      RECT 65.145 72.417 65.211 74.722 ;
      RECT 62.937 74.625 65.257 74.676 ;
      RECT 65.191 72.371 65.257 74.676 ;
      RECT 62.983 74.579 65.303 74.63 ;
      RECT 65.237 72.325 65.303 74.63 ;
      RECT 63.029 74.533 65.349 74.584 ;
      RECT 65.283 72.279 65.349 74.584 ;
      RECT 63.075 74.487 65.395 74.538 ;
      RECT 65.329 72.233 65.395 74.538 ;
      RECT 63.121 74.441 65.441 74.492 ;
      RECT 65.375 72.187 65.441 74.492 ;
      RECT 63.167 74.395 65.487 74.446 ;
      RECT 65.421 72.141 65.487 74.446 ;
      RECT 63.213 74.349 65.533 74.4 ;
      RECT 65.467 72.095 65.533 74.4 ;
      RECT 63.259 74.303 65.579 74.354 ;
      RECT 65.513 72.049 65.579 74.354 ;
      RECT 65.559 72.003 65.625 74.308 ;
      RECT 65.605 71.957 65.671 74.262 ;
      RECT 65.651 71.911 65.717 74.216 ;
      RECT 65.697 71.865 65.763 74.17 ;
      RECT 65.743 71.819 65.809 74.124 ;
      RECT 65.789 71.773 65.855 74.078 ;
      RECT 65.835 71.727 65.901 74.032 ;
      RECT 65.881 71.681 65.947 73.986 ;
      RECT 65.927 71.635 65.993 73.94 ;
      RECT 65.973 71.589 66.039 73.894 ;
      RECT 66.019 71.543 66.085 73.848 ;
      RECT 66.065 71.497 66.131 73.802 ;
      RECT 66.111 71.451 66.177 73.756 ;
      RECT 66.157 71.405 66.223 73.71 ;
      RECT 66.203 71.359 66.269 73.664 ;
      RECT 66.249 71.313 66.315 73.618 ;
      RECT 66.295 71.267 66.361 73.572 ;
      RECT 66.341 71.221 66.407 73.526 ;
      RECT 66.387 71.175 66.453 73.48 ;
      RECT 66.433 71.129 66.499 73.434 ;
      RECT 66.479 71.083 66.545 73.388 ;
      RECT 66.525 71.037 66.591 73.342 ;
      RECT 66.571 70.991 66.637 73.296 ;
      RECT 66.617 70.945 66.683 73.25 ;
      RECT 66.663 70.899 66.729 73.204 ;
      RECT 66.709 70.853 66.775 73.158 ;
      RECT 66.755 70.807 66.821 73.112 ;
      RECT 66.801 70.761 66.867 73.066 ;
      RECT 66.847 70.715 66.913 73.02 ;
      RECT 66.893 70.669 66.959 72.974 ;
      RECT 66.939 70.623 67.005 72.928 ;
      RECT 66.985 70.577 67.051 72.882 ;
      RECT 67.031 70.531 67.097 72.836 ;
      RECT 67.077 70.485 67.143 72.79 ;
      RECT 67.123 70.439 67.189 72.744 ;
      RECT 67.169 70.393 67.235 72.698 ;
      RECT 67.215 70.347 67.281 72.652 ;
      RECT 67.261 70.301 67.327 72.606 ;
      RECT 67.307 70.255 67.373 72.56 ;
      RECT 67.353 70.209 67.419 72.514 ;
      RECT 67.399 70.163 67.465 72.468 ;
      RECT 67.445 70.117 67.511 72.422 ;
      RECT 67.491 70.071 67.557 72.376 ;
      RECT 67.537 70.025 67.603 72.33 ;
      RECT 67.583 69.979 67.649 72.284 ;
      RECT 67.629 69.933 67.695 72.238 ;
      RECT 67.675 69.887 67.741 72.192 ;
      RECT 67.721 69.841 67.787 72.146 ;
      RECT 67.767 69.795 67.833 72.1 ;
      RECT 67.813 69.749 67.879 72.054 ;
      RECT 67.859 69.703 67.925 72.008 ;
      RECT 67.905 69.657 67.971 71.962 ;
      RECT 67.951 69.611 68.017 71.916 ;
      RECT 67.997 69.565 68.063 71.87 ;
      RECT 68.043 69.519 68.109 71.824 ;
      RECT 68.089 69.473 68.155 71.778 ;
      RECT 68.135 69.427 68.201 71.732 ;
      RECT 68.181 69.381 68.247 71.686 ;
      RECT 68.227 69.335 68.293 71.64 ;
      RECT 68.273 69.289 68.339 71.594 ;
      RECT 68.319 69.243 68.385 71.548 ;
      RECT 68.365 69.197 68.431 71.502 ;
      RECT 68.411 69.151 68.477 71.456 ;
      RECT 68.457 69.105 68.523 71.41 ;
      RECT 68.503 69.059 68.569 71.364 ;
      RECT 68.549 69.013 68.615 71.318 ;
      RECT 68.595 68.967 68.661 71.272 ;
      RECT 68.641 68.921 68.707 71.226 ;
      RECT 68.687 68.875 68.753 71.18 ;
      RECT 68.733 68.829 68.799 71.134 ;
      RECT 68.779 68.783 68.845 71.088 ;
      RECT 68.825 68.737 68.891 71.042 ;
      RECT 68.871 68.691 68.937 70.996 ;
      RECT 68.917 68.645 68.983 70.95 ;
      RECT 68.963 68.599 69.029 70.904 ;
      RECT 69.009 68.553 69.075 70.858 ;
      RECT 69.055 68.507 69.121 70.812 ;
      RECT 69.101 68.461 69.167 70.766 ;
      RECT 69.147 68.415 69.213 70.72 ;
      RECT 69.193 68.369 69.259 70.674 ;
      RECT 69.239 68.323 69.305 70.628 ;
      RECT 69.285 68.277 69.351 70.582 ;
      RECT 69.331 68.231 69.397 70.536 ;
      RECT 69.377 68.185 69.443 70.49 ;
      RECT 69.423 68.139 69.489 70.444 ;
      RECT 69.469 68.093 69.535 70.398 ;
      RECT 69.515 68.047 69.581 70.352 ;
      RECT 69.561 68.001 69.627 70.306 ;
      RECT 69.607 67.955 69.673 70.26 ;
      RECT 69.653 67.909 69.719 70.214 ;
      RECT 69.699 67.863 69.765 70.168 ;
      RECT 69.745 67.817 69.811 70.122 ;
      RECT 69.791 67.771 69.857 70.076 ;
      RECT 69.837 67.725 69.903 70.03 ;
      RECT 69.883 67.679 69.949 69.984 ;
      RECT 69.929 67.633 69.995 69.938 ;
      RECT 69.975 67.587 70.041 69.892 ;
      RECT 70.021 67.541 70.087 69.846 ;
      RECT 70.067 67.495 70.133 69.8 ;
      RECT 70.113 67.449 70.179 69.754 ;
      RECT 70.159 67.403 70.225 69.708 ;
      RECT 70.205 67.357 70.271 69.662 ;
      RECT 70.251 67.311 70.317 69.616 ;
      RECT 70.297 67.265 70.363 69.57 ;
      RECT 70.343 67.219 70.409 69.524 ;
      RECT 70.389 67.173 70.455 69.478 ;
      RECT 70.435 67.127 70.501 69.432 ;
      RECT 70.481 67.081 70.547 69.386 ;
      RECT 70.527 67.035 70.593 69.34 ;
      RECT 70.573 66.989 70.639 69.294 ;
      RECT 70.619 66.943 70.685 69.248 ;
      RECT 70.665 66.897 70.731 69.202 ;
      RECT 70.711 66.851 70.777 69.156 ;
      RECT 70.757 66.805 70.823 69.11 ;
      RECT 70.803 66.759 70.869 69.064 ;
      RECT 70.849 66.713 70.915 69.018 ;
      RECT 70.895 66.667 70.961 68.972 ;
      RECT 70.941 66.621 71.007 68.926 ;
      RECT 70.987 66.575 71.053 68.88 ;
      RECT 71.033 66.529 71.099 68.834 ;
      RECT 71.079 66.483 71.145 68.788 ;
      RECT 71.125 66.437 71.191 68.742 ;
      RECT 71.171 66.391 71.237 68.696 ;
      RECT 71.217 66.345 71.283 68.65 ;
      RECT 71.263 66.299 71.329 68.604 ;
      RECT 71.309 66.253 71.375 68.558 ;
      RECT 71.355 66.207 71.421 68.512 ;
      RECT 71.401 66.161 71.467 68.466 ;
      RECT 71.447 66.115 71.513 68.42 ;
      RECT 71.493 66.069 71.559 68.374 ;
      RECT 71.539 66.023 71.605 68.328 ;
      RECT 71.585 65.977 71.651 68.282 ;
      RECT 71.631 65.931 71.697 68.236 ;
      RECT 71.677 65.885 71.743 68.19 ;
      RECT 71.723 65.839 71.789 68.144 ;
      RECT 71.769 65.793 71.835 68.098 ;
      RECT 71.815 65.747 71.881 68.052 ;
      RECT 71.861 65.701 71.927 68.006 ;
      RECT 71.907 65.655 71.973 67.96 ;
      RECT 71.953 65.609 72.019 67.914 ;
      RECT 71.999 65.563 72.065 67.868 ;
      RECT 72.045 65.517 72.111 67.822 ;
      RECT 72.091 65.471 72.157 67.776 ;
      RECT 72.137 65.425 72.203 67.73 ;
      RECT 72.183 65.379 72.249 67.684 ;
      RECT 72.229 65.333 72.295 67.638 ;
      RECT 72.275 65.287 72.341 67.592 ;
      RECT 72.321 65.241 72.387 67.546 ;
      RECT 72.367 65.195 72.433 67.5 ;
      RECT 72.413 65.149 72.479 67.454 ;
      RECT 72.459 65.103 72.525 67.408 ;
      RECT 72.505 65.057 72.571 67.362 ;
      RECT 72.551 65.011 72.617 67.316 ;
      RECT 72.597 64.965 72.663 67.27 ;
      RECT 72.643 64.919 72.709 67.224 ;
      RECT 72.689 64.873 72.755 67.178 ;
      RECT 72.735 64.827 72.801 67.132 ;
      RECT 72.781 64.781 72.847 67.086 ;
      RECT 72.827 64.735 72.893 67.04 ;
      RECT 72.873 64.689 72.939 66.994 ;
      RECT 72.919 64.643 72.985 66.948 ;
      RECT 72.965 64.597 73.031 66.902 ;
      RECT 73.011 64.551 73.077 66.856 ;
      RECT 73.057 64.505 73.123 66.81 ;
      RECT 73.103 64.459 73.169 66.764 ;
      RECT 73.149 64.413 73.215 66.718 ;
      RECT 73.195 64.367 73.261 66.672 ;
      RECT 73.241 64.321 73.307 66.626 ;
      RECT 73.287 64.275 73.353 66.58 ;
      RECT 73.333 64.229 73.399 66.534 ;
      RECT 73.379 64.183 73.445 66.488 ;
      RECT 73.425 64.137 73.491 66.442 ;
      RECT 73.471 64.091 73.537 66.396 ;
      RECT 73.517 64.045 73.583 66.35 ;
      RECT 73.563 63.999 73.629 66.304 ;
      RECT 73.609 63.953 73.675 66.258 ;
      RECT 73.655 63.907 73.721 66.212 ;
      RECT 73.701 63.861 73.767 66.166 ;
      RECT 73.747 63.815 73.813 66.12 ;
      RECT 73.793 63.769 73.859 66.074 ;
      RECT 73.839 63.723 73.905 66.028 ;
      RECT 73.885 63.677 73.951 65.982 ;
      RECT 73.931 63.631 73.997 65.936 ;
      RECT 73.977 63.585 74.043 65.89 ;
      RECT 74.023 63.539 74.089 65.844 ;
      RECT 74.069 63.493 74.135 65.798 ;
      RECT 74.115 63.447 74.181 65.752 ;
      RECT 74.161 63.401 74.227 65.706 ;
      RECT 74.207 63.355 74.273 65.66 ;
      RECT 74.253 63.309 74.319 65.614 ;
      RECT 74.299 63.263 74.365 65.568 ;
      RECT 74.345 63.217 74.411 65.522 ;
      RECT 74.391 63.171 74.457 65.476 ;
      RECT 74.437 63.125 74.503 65.43 ;
      RECT 74.483 63.079 74.549 65.384 ;
      RECT 74.529 63.033 74.595 65.338 ;
      RECT 74.575 62.987 74.641 65.292 ;
      RECT 74.621 62.941 74.687 65.246 ;
      RECT 74.667 62.895 74.733 65.2 ;
      RECT 74.713 62.849 74.779 65.154 ;
      RECT 74.759 62.803 74.825 65.108 ;
      RECT 74.805 62.757 74.871 65.062 ;
      RECT 74.851 62.711 74.917 65.016 ;
      RECT 74.897 62.665 74.963 64.97 ;
      RECT 74.943 62.619 75.009 64.924 ;
      RECT 74.989 62.573 75.055 64.878 ;
      RECT 75.035 62.527 75.101 64.832 ;
      RECT 75.081 62.481 75.147 64.786 ;
      RECT 75.127 62.435 75.193 64.74 ;
      RECT 75.173 62.389 75.239 64.694 ;
      RECT 75.219 62.343 75.285 64.648 ;
      RECT 75.265 62.297 75.331 64.602 ;
      RECT 75.311 62.251 75.377 64.556 ;
      RECT 75.357 62.205 75.423 64.51 ;
      RECT 75.403 62.159 75.469 64.464 ;
      RECT 75.449 62.113 75.515 64.418 ;
      RECT 75.495 62.067 75.561 64.372 ;
      RECT 75.541 62.021 75.607 64.326 ;
      RECT 75.587 61.975 75.653 64.28 ;
      RECT 75.633 61.929 75.699 64.234 ;
      RECT 75.679 61.883 75.745 64.188 ;
      RECT 75.725 61.837 75.791 64.142 ;
      RECT 75.771 61.791 75.837 64.096 ;
      RECT 75.817 61.745 75.883 64.05 ;
      RECT 75.863 61.699 75.929 64.004 ;
      RECT 75.909 61.653 75.975 63.958 ;
      RECT 75.955 61.607 76.021 63.912 ;
      RECT 76.001 61.561 76.067 63.866 ;
      RECT 76.047 61.515 76.113 63.82 ;
      RECT 76.093 61.469 76.159 63.774 ;
      RECT 76.139 61.423 76.205 63.728 ;
      RECT 76.185 61.377 76.251 63.682 ;
      RECT 76.231 61.331 76.297 63.636 ;
      RECT 76.277 61.285 76.343 63.59 ;
      RECT 76.323 61.239 76.389 63.544 ;
      RECT 76.369 61.193 76.435 63.498 ;
      RECT 76.415 61.158 76.481 63.452 ;
      RECT 76.44 61.122 76.527 63.406 ;
      RECT 76.486 61.076 76.573 63.36 ;
      RECT 76.532 61.03 76.619 63.314 ;
      RECT 76.578 60.984 76.665 63.268 ;
      RECT 76.624 60.938 76.711 63.222 ;
      RECT 76.67 60.892 76.757 63.176 ;
      RECT 76.716 60.846 76.803 63.13 ;
      RECT 76.762 60.8 76.849 63.084 ;
      RECT 76.808 60.754 76.895 63.038 ;
      RECT 76.854 60.708 76.941 62.992 ;
      RECT 76.9 60.662 76.987 62.946 ;
      RECT 76.946 60.616 77.033 62.9 ;
      RECT 76.992 60.57 77.079 62.854 ;
      RECT 77.038 60.524 77.125 62.808 ;
      RECT 77.084 60.478 77.171 62.762 ;
      RECT 77.13 60.432 77.217 62.716 ;
      RECT 77.176 60.386 77.263 62.67 ;
      RECT 77.222 60.34 77.309 62.624 ;
      RECT 77.268 60.294 77.355 62.578 ;
      RECT 77.314 60.248 77.401 62.532 ;
      RECT 77.36 60.202 77.447 62.486 ;
      RECT 77.406 60.156 77.493 62.44 ;
      RECT 77.452 60.11 77.539 62.394 ;
      RECT 77.498 60.064 77.585 62.348 ;
      RECT 77.544 60.018 77.631 62.302 ;
      RECT 77.59 59.972 77.677 62.256 ;
      RECT 77.636 59.926 77.723 62.21 ;
      RECT 77.682 59.88 77.769 62.164 ;
      RECT 77.728 59.834 77.815 62.118 ;
      RECT 77.774 59.788 77.861 62.072 ;
      RECT 77.82 59.742 77.907 62.026 ;
      RECT 77.866 59.696 77.953 61.98 ;
      RECT 77.912 59.65 77.999 61.934 ;
      RECT 77.958 59.604 78.045 61.888 ;
      RECT 78.004 59.558 78.091 61.842 ;
      RECT 78.05 59.512 78.137 61.796 ;
      RECT 78.096 59.466 78.183 61.75 ;
      RECT 78.142 59.42 78.229 61.704 ;
      RECT 78.188 59.374 78.275 61.658 ;
      RECT 78.234 59.328 78.321 61.612 ;
      RECT 78.28 59.282 78.367 61.566 ;
      RECT 78.326 59.236 78.413 61.52 ;
      RECT 78.372 59.19 78.459 61.474 ;
      RECT 78.418 59.144 78.505 61.428 ;
      RECT 78.464 59.098 78.551 61.382 ;
      RECT 78.51 59.052 78.597 61.336 ;
      RECT 78.556 59.006 78.643 61.29 ;
      RECT 78.602 58.96 78.689 61.244 ;
      RECT 78.648 58.914 78.735 61.198 ;
      RECT 78.694 58.868 78.781 61.152 ;
      RECT 78.74 58.822 78.827 61.106 ;
      RECT 78.786 58.776 78.873 61.06 ;
      RECT 78.832 58.73 78.919 61.014 ;
      RECT 78.878 58.684 78.965 60.968 ;
      RECT 78.924 58.638 79.011 60.922 ;
      RECT 78.97 58.592 79.057 60.876 ;
      RECT 79.016 58.546 79.103 60.83 ;
      RECT 79.062 58.5 79.149 60.784 ;
      RECT 79.108 58.454 79.195 60.738 ;
      RECT 79.154 58.408 79.241 60.692 ;
      RECT 79.2 58.362 79.287 60.646 ;
      RECT 79.246 58.316 79.333 60.6 ;
      RECT 79.292 58.27 79.379 60.554 ;
      RECT 79.338 58.224 79.425 60.508 ;
      RECT 79.384 58.178 79.471 60.462 ;
      RECT 79.43 58.132 79.517 60.416 ;
      RECT 79.476 58.086 79.563 60.37 ;
      RECT 79.522 58.04 79.609 60.324 ;
      RECT 79.568 57.994 79.655 60.278 ;
      RECT 79.614 57.948 79.701 60.232 ;
      RECT 79.66 57.902 79.747 60.186 ;
      RECT 79.706 57.856 79.793 60.14 ;
      RECT 79.752 57.81 79.839 60.094 ;
      RECT 79.798 57.764 79.885 60.048 ;
      RECT 79.844 57.718 79.931 60.002 ;
      RECT 79.89 57.672 79.977 59.956 ;
      RECT 79.936 57.626 80.023 59.91 ;
      RECT 79.982 57.58 80.069 59.864 ;
      RECT 80.028 57.534 80.115 59.818 ;
      RECT 80.074 57.488 80.161 59.772 ;
      RECT 80.12 57.442 80.207 59.726 ;
      RECT 80.166 57.396 80.253 59.68 ;
      RECT 80.212 57.35 80.299 59.634 ;
      RECT 80.258 57.304 80.345 59.588 ;
      RECT 80.304 57.258 80.391 59.542 ;
      RECT 80.35 57.212 80.437 59.496 ;
      RECT 80.396 57.166 80.483 59.45 ;
      RECT 80.442 57.12 80.529 59.404 ;
      RECT 80.488 57.074 80.575 59.358 ;
      RECT 80.534 57.028 80.621 59.312 ;
      RECT 80.58 56.982 80.667 59.266 ;
      RECT 80.626 56.936 80.713 59.22 ;
      RECT 80.672 56.89 80.759 59.174 ;
      RECT 80.718 56.844 80.805 59.128 ;
      RECT 80.764 56.798 80.851 59.082 ;
      RECT 80.81 56.752 80.897 59.036 ;
      RECT 80.856 56.706 80.943 58.99 ;
      RECT 80.902 56.66 80.989 58.944 ;
      RECT 80.948 56.614 81.035 58.898 ;
      RECT 80.994 56.568 81.081 58.852 ;
      RECT 81.04 56.522 81.127 58.806 ;
      RECT 81.086 56.476 81.173 58.76 ;
      RECT 81.132 56.43 81.219 58.714 ;
      RECT 81.178 56.384 81.265 58.668 ;
      RECT 81.224 56.338 81.311 58.622 ;
      RECT 81.27 56.292 81.357 58.576 ;
      RECT 81.316 56.246 81.403 58.53 ;
      RECT 81.362 56.199 81.449 58.484 ;
      RECT 81.408 56.175 81.495 58.438 ;
      RECT 81.408 56.175 81.541 58.392 ;
      RECT 81.408 56.175 81.587 58.346 ;
      RECT 81.408 56.175 81.633 58.3 ;
      RECT 81.408 56.175 81.679 58.254 ;
      RECT 81.408 56.175 81.725 58.208 ;
      RECT 81.408 56.175 81.771 58.162 ;
      RECT 81.408 56.175 81.817 58.116 ;
      RECT 81.408 56.175 81.863 58.07 ;
      RECT 81.408 56.175 81.909 58.024 ;
      RECT 81.408 56.175 81.955 57.978 ;
      RECT 81.408 56.175 82.001 57.932 ;
      RECT 81.408 56.175 82.047 57.886 ;
      RECT 81.408 56.175 82.093 57.84 ;
      RECT 81.408 56.175 82.139 57.794 ;
      RECT 81.408 56.175 82.185 57.748 ;
      RECT 81.408 56.175 82.231 57.702 ;
      RECT 81.408 56.175 82.277 57.656 ;
      RECT 81.408 56.175 82.323 57.61 ;
      RECT 81.408 56.175 82.369 57.564 ;
      RECT 81.408 56.175 82.415 57.518 ;
      RECT 81.408 56.175 82.461 57.472 ;
      RECT 81.408 56.175 82.507 57.426 ;
      RECT 81.408 56.175 82.553 57.38 ;
      RECT 80.258 57.304 82.585 57.341 ;
      RECT 81.408 56.175 110 57.325 ;
      RECT 63.675 85.392 68.325 110 ;
      RECT 63.675 85.392 68.371 88.167 ;
      RECT 63.675 85.392 68.417 88.121 ;
      RECT 63.675 85.392 68.463 88.075 ;
      RECT 63.675 85.392 68.509 88.029 ;
      RECT 63.675 85.392 68.555 87.983 ;
      RECT 63.675 85.392 68.601 87.937 ;
      RECT 63.675 85.392 68.647 87.891 ;
      RECT 63.675 85.392 68.693 87.845 ;
      RECT 63.675 85.392 68.739 87.799 ;
      RECT 63.675 85.392 68.785 87.753 ;
      RECT 63.675 85.392 68.831 87.707 ;
      RECT 63.675 85.392 68.877 87.661 ;
      RECT 63.675 85.392 68.923 87.615 ;
      RECT 63.675 85.392 68.969 87.569 ;
      RECT 63.675 85.392 69.015 87.523 ;
      RECT 63.675 85.392 69.061 87.477 ;
      RECT 63.675 85.392 69.107 87.431 ;
      RECT 63.675 85.392 69.153 87.385 ;
      RECT 63.675 85.392 69.199 87.339 ;
      RECT 63.675 85.392 69.245 87.293 ;
      RECT 63.675 85.392 69.291 87.247 ;
      RECT 63.675 85.392 69.337 87.201 ;
      RECT 63.675 85.392 69.383 87.155 ;
      RECT 63.675 85.392 69.429 87.109 ;
      RECT 63.675 85.392 69.475 87.063 ;
      RECT 63.675 85.392 69.521 87.017 ;
      RECT 63.675 85.392 69.567 86.971 ;
      RECT 63.675 85.392 69.613 86.925 ;
      RECT 63.675 85.392 69.659 86.879 ;
      RECT 63.675 85.392 69.705 86.833 ;
      RECT 63.675 85.392 69.751 86.787 ;
      RECT 63.675 85.392 69.797 86.741 ;
      RECT 63.675 85.392 69.843 86.695 ;
      RECT 63.675 85.392 69.889 86.649 ;
      RECT 63.675 85.392 69.935 86.603 ;
      RECT 63.675 85.392 69.981 86.557 ;
      RECT 63.675 85.392 70.027 86.511 ;
      RECT 63.675 85.392 70.073 86.465 ;
      RECT 63.675 85.392 70.119 86.419 ;
      RECT 63.675 85.392 70.165 86.373 ;
      RECT 63.675 85.392 70.211 86.327 ;
      RECT 63.675 85.392 70.257 86.281 ;
      RECT 63.675 85.392 70.303 86.235 ;
      RECT 63.675 85.392 70.349 86.189 ;
      RECT 63.675 85.392 70.395 86.143 ;
      RECT 63.675 85.392 70.441 86.097 ;
      RECT 63.675 85.392 70.487 86.051 ;
      RECT 63.675 85.392 70.533 86.005 ;
      RECT 63.675 85.392 70.579 85.959 ;
      RECT 63.675 85.392 70.625 85.913 ;
      RECT 63.675 85.392 70.671 85.867 ;
      RECT 63.675 85.392 70.717 85.821 ;
      RECT 63.675 85.392 70.763 85.775 ;
      RECT 63.675 85.392 70.809 85.729 ;
      RECT 63.675 85.392 70.855 85.683 ;
      RECT 63.675 85.392 70.901 85.637 ;
      RECT 63.675 85.392 70.947 85.591 ;
      RECT 63.675 85.392 70.993 85.545 ;
      RECT 63.675 85.392 71.039 85.499 ;
      RECT 63.721 85.346 71.131 85.407 ;
      RECT 71.081 77.986 71.131 85.407 ;
      RECT 63.767 85.3 71.177 85.361 ;
      RECT 71.127 77.94 71.177 85.361 ;
      RECT 63.813 85.254 71.223 85.315 ;
      RECT 71.173 77.894 71.223 85.315 ;
      RECT 63.859 85.208 71.269 85.269 ;
      RECT 71.219 77.848 71.269 85.269 ;
      RECT 63.905 85.162 71.315 85.223 ;
      RECT 71.265 77.802 71.315 85.223 ;
      RECT 63.951 85.116 71.361 85.177 ;
      RECT 71.311 77.756 71.361 85.177 ;
      RECT 63.997 85.07 71.407 85.131 ;
      RECT 71.357 77.71 71.407 85.131 ;
      RECT 64.043 85.024 71.453 85.085 ;
      RECT 71.403 77.664 71.453 85.085 ;
      RECT 64.089 84.978 71.499 85.039 ;
      RECT 71.449 77.618 71.499 85.039 ;
      RECT 64.135 84.932 71.545 84.993 ;
      RECT 71.495 77.572 71.545 84.993 ;
      RECT 64.181 84.886 71.591 84.947 ;
      RECT 71.541 77.526 71.591 84.947 ;
      RECT 64.227 84.84 71.637 84.901 ;
      RECT 71.587 77.48 71.637 84.901 ;
      RECT 64.273 84.794 71.683 84.855 ;
      RECT 71.633 77.434 71.683 84.855 ;
      RECT 64.319 84.748 71.729 84.809 ;
      RECT 71.679 77.388 71.729 84.809 ;
      RECT 64.365 84.702 71.775 84.763 ;
      RECT 71.725 77.342 71.775 84.763 ;
      RECT 64.411 84.656 71.821 84.717 ;
      RECT 71.771 77.296 71.821 84.717 ;
      RECT 64.457 84.61 71.867 84.671 ;
      RECT 71.817 77.25 71.867 84.671 ;
      RECT 64.503 84.564 71.913 84.625 ;
      RECT 71.863 77.204 71.913 84.625 ;
      RECT 64.549 84.518 71.959 84.579 ;
      RECT 71.909 77.158 71.959 84.579 ;
      RECT 64.595 84.472 72.005 84.533 ;
      RECT 71.955 77.112 72.005 84.533 ;
      RECT 64.641 84.426 72.051 84.487 ;
      RECT 72.001 77.066 72.051 84.487 ;
      RECT 64.687 84.38 72.097 84.441 ;
      RECT 72.047 77.02 72.097 84.441 ;
      RECT 64.733 84.334 72.143 84.395 ;
      RECT 72.093 76.974 72.143 84.395 ;
      RECT 64.779 84.288 72.189 84.349 ;
      RECT 72.139 76.928 72.189 84.349 ;
      RECT 64.825 84.242 72.235 84.303 ;
      RECT 72.185 76.882 72.235 84.303 ;
      RECT 64.871 84.196 72.281 84.257 ;
      RECT 72.231 76.836 72.281 84.257 ;
      RECT 64.917 84.15 72.327 84.211 ;
      RECT 72.277 76.79 72.327 84.211 ;
      RECT 64.963 84.104 72.373 84.165 ;
      RECT 72.323 76.744 72.373 84.165 ;
      RECT 65.009 84.058 72.419 84.119 ;
      RECT 72.369 76.698 72.419 84.119 ;
      RECT 65.055 84.012 72.465 84.073 ;
      RECT 72.415 76.652 72.465 84.073 ;
      RECT 65.101 83.966 72.511 84.027 ;
      RECT 72.461 76.606 72.511 84.027 ;
      RECT 65.147 83.92 72.557 83.981 ;
      RECT 72.507 76.56 72.557 83.981 ;
      RECT 65.193 83.874 72.603 83.935 ;
      RECT 72.553 76.514 72.603 83.935 ;
      RECT 65.239 83.828 72.649 83.889 ;
      RECT 72.599 76.468 72.649 83.889 ;
      RECT 65.285 83.782 72.695 83.843 ;
      RECT 72.645 76.422 72.695 83.843 ;
      RECT 65.331 83.736 72.741 83.797 ;
      RECT 72.691 76.376 72.741 83.797 ;
      RECT 65.377 83.69 72.787 83.751 ;
      RECT 72.737 76.33 72.787 83.751 ;
      RECT 65.423 83.644 72.833 83.705 ;
      RECT 72.783 76.284 72.833 83.705 ;
      RECT 65.469 83.598 72.879 83.659 ;
      RECT 72.829 76.238 72.879 83.659 ;
      RECT 65.515 83.552 72.925 83.613 ;
      RECT 72.875 76.192 72.925 83.613 ;
      RECT 65.561 83.506 72.971 83.567 ;
      RECT 72.921 76.146 72.971 83.567 ;
      RECT 65.607 83.46 73.017 83.521 ;
      RECT 72.967 76.1 73.017 83.521 ;
      RECT 65.653 83.414 73.063 83.475 ;
      RECT 73.013 76.054 73.063 83.475 ;
      RECT 65.699 83.368 73.109 83.429 ;
      RECT 73.059 76.008 73.109 83.429 ;
      RECT 65.745 83.322 73.155 83.383 ;
      RECT 73.105 75.962 73.155 83.383 ;
      RECT 65.791 83.276 73.201 83.337 ;
      RECT 73.151 75.916 73.201 83.337 ;
      RECT 65.837 83.23 73.247 83.291 ;
      RECT 73.197 75.87 73.247 83.291 ;
      RECT 65.883 83.184 73.293 83.245 ;
      RECT 73.243 75.824 73.293 83.245 ;
      RECT 65.929 83.138 73.339 83.199 ;
      RECT 73.289 75.778 73.339 83.199 ;
      RECT 65.975 83.092 73.385 83.153 ;
      RECT 73.335 75.732 73.385 83.153 ;
      RECT 66.021 83.046 73.431 83.107 ;
      RECT 73.381 75.686 73.431 83.107 ;
      RECT 66.067 83 73.477 83.061 ;
      RECT 73.427 75.64 73.477 83.061 ;
      RECT 66.113 82.954 73.523 83.015 ;
      RECT 73.473 75.594 73.523 83.015 ;
      RECT 66.159 82.908 73.569 82.969 ;
      RECT 73.519 75.548 73.569 82.969 ;
      RECT 66.205 82.862 73.615 82.923 ;
      RECT 73.565 75.502 73.615 82.923 ;
      RECT 66.251 82.816 73.661 82.877 ;
      RECT 73.611 75.456 73.661 82.877 ;
      RECT 66.297 82.77 73.707 82.831 ;
      RECT 73.657 75.41 73.707 82.831 ;
      RECT 66.343 82.724 73.753 82.785 ;
      RECT 73.703 75.364 73.753 82.785 ;
      RECT 66.389 82.678 73.799 82.739 ;
      RECT 73.749 75.318 73.799 82.739 ;
      RECT 66.435 82.632 73.845 82.693 ;
      RECT 73.795 75.272 73.845 82.693 ;
      RECT 66.481 82.586 73.891 82.647 ;
      RECT 73.841 75.226 73.891 82.647 ;
      RECT 66.527 82.54 73.937 82.601 ;
      RECT 73.887 75.18 73.937 82.601 ;
      RECT 66.573 82.494 73.983 82.555 ;
      RECT 73.933 75.134 73.983 82.555 ;
      RECT 66.619 82.448 74.029 82.509 ;
      RECT 73.979 75.088 74.029 82.509 ;
      RECT 66.665 82.402 74.075 82.463 ;
      RECT 74.025 75.042 74.075 82.463 ;
      RECT 66.711 82.356 74.121 82.417 ;
      RECT 74.071 74.996 74.121 82.417 ;
      RECT 66.757 82.31 74.167 82.371 ;
      RECT 74.117 74.95 74.167 82.371 ;
      RECT 66.803 82.264 74.213 82.325 ;
      RECT 74.163 74.904 74.213 82.325 ;
      RECT 66.849 82.218 74.259 82.279 ;
      RECT 74.209 74.858 74.259 82.279 ;
      RECT 66.895 82.172 74.305 82.233 ;
      RECT 74.255 74.812 74.305 82.233 ;
      RECT 66.941 82.126 74.351 82.187 ;
      RECT 74.301 74.766 74.351 82.187 ;
      RECT 66.987 82.08 74.397 82.141 ;
      RECT 74.347 74.72 74.397 82.141 ;
      RECT 67.033 82.034 74.443 82.095 ;
      RECT 74.393 74.674 74.443 82.095 ;
      RECT 67.079 81.988 74.489 82.049 ;
      RECT 74.439 74.628 74.489 82.049 ;
      RECT 67.125 81.942 74.535 82.003 ;
      RECT 74.485 74.582 74.535 82.003 ;
      RECT 67.171 81.896 74.581 81.957 ;
      RECT 74.531 74.536 74.581 81.957 ;
      RECT 67.217 81.85 74.627 81.911 ;
      RECT 74.577 74.49 74.627 81.911 ;
      RECT 67.263 81.804 74.673 81.865 ;
      RECT 74.623 74.444 74.673 81.865 ;
      RECT 67.309 81.758 74.719 81.819 ;
      RECT 74.669 74.398 74.719 81.819 ;
      RECT 67.355 81.712 74.765 81.773 ;
      RECT 74.715 74.352 74.765 81.773 ;
      RECT 67.401 81.666 74.811 81.727 ;
      RECT 74.761 74.306 74.811 81.727 ;
      RECT 67.447 81.62 74.857 81.681 ;
      RECT 74.807 74.26 74.857 81.681 ;
      RECT 67.493 81.574 74.903 81.635 ;
      RECT 74.853 74.214 74.903 81.635 ;
      RECT 67.539 81.528 74.949 81.589 ;
      RECT 74.899 74.168 74.949 81.589 ;
      RECT 67.585 81.482 74.995 81.543 ;
      RECT 74.945 74.122 74.995 81.543 ;
      RECT 67.631 81.436 75.041 81.497 ;
      RECT 74.991 74.076 75.041 81.497 ;
      RECT 67.677 81.39 75.087 81.451 ;
      RECT 75.037 74.03 75.087 81.451 ;
      RECT 67.723 81.344 75.133 81.405 ;
      RECT 75.083 73.984 75.133 81.405 ;
      RECT 67.769 81.298 75.179 81.359 ;
      RECT 75.129 73.938 75.179 81.359 ;
      RECT 67.815 81.252 75.225 81.313 ;
      RECT 75.175 73.892 75.225 81.313 ;
      RECT 67.861 81.206 75.271 81.267 ;
      RECT 75.221 73.846 75.271 81.267 ;
      RECT 67.907 81.16 75.317 81.221 ;
      RECT 75.267 73.8 75.317 81.221 ;
      RECT 67.953 81.114 75.363 81.175 ;
      RECT 75.313 73.754 75.363 81.175 ;
      RECT 67.999 81.068 75.409 81.129 ;
      RECT 75.359 73.708 75.409 81.129 ;
      RECT 68.045 81.022 75.455 81.083 ;
      RECT 75.405 73.662 75.455 81.083 ;
      RECT 68.091 80.976 75.501 81.037 ;
      RECT 75.451 73.616 75.501 81.037 ;
      RECT 68.137 80.93 75.547 80.991 ;
      RECT 75.497 73.57 75.547 80.991 ;
      RECT 68.183 80.884 75.593 80.945 ;
      RECT 75.543 73.524 75.593 80.945 ;
      RECT 68.229 80.838 75.639 80.899 ;
      RECT 75.589 73.478 75.639 80.899 ;
      RECT 68.275 80.792 75.685 80.853 ;
      RECT 75.635 73.432 75.685 80.853 ;
      RECT 68.321 80.746 75.731 80.807 ;
      RECT 75.681 73.386 75.731 80.807 ;
      RECT 68.367 80.7 75.777 80.761 ;
      RECT 75.727 73.34 75.777 80.761 ;
      RECT 68.413 80.654 75.823 80.715 ;
      RECT 75.773 73.294 75.823 80.715 ;
      RECT 68.459 80.608 75.869 80.669 ;
      RECT 75.819 73.248 75.869 80.669 ;
      RECT 68.505 80.562 75.915 80.623 ;
      RECT 75.865 73.202 75.915 80.623 ;
      RECT 68.551 80.516 75.961 80.577 ;
      RECT 75.911 73.156 75.961 80.577 ;
      RECT 68.597 80.47 76.007 80.531 ;
      RECT 75.957 73.11 76.007 80.531 ;
      RECT 68.643 80.424 76.053 80.485 ;
      RECT 76.003 73.064 76.053 80.485 ;
      RECT 68.689 80.378 76.099 80.439 ;
      RECT 76.049 73.018 76.099 80.439 ;
      RECT 68.735 80.332 76.145 80.393 ;
      RECT 76.095 72.972 76.145 80.393 ;
      RECT 68.781 80.286 76.191 80.347 ;
      RECT 76.141 72.926 76.191 80.347 ;
      RECT 68.827 80.24 76.237 80.301 ;
      RECT 76.187 72.88 76.237 80.301 ;
      RECT 68.873 80.194 76.283 80.255 ;
      RECT 76.233 72.834 76.283 80.255 ;
      RECT 68.919 80.148 76.329 80.209 ;
      RECT 76.279 72.788 76.329 80.209 ;
      RECT 68.965 80.102 76.375 80.163 ;
      RECT 76.325 72.742 76.375 80.163 ;
      RECT 69.011 80.056 76.421 80.117 ;
      RECT 76.371 72.696 76.421 80.117 ;
      RECT 69.057 80.01 76.467 80.071 ;
      RECT 76.417 72.65 76.467 80.071 ;
      RECT 69.103 79.964 76.513 80.025 ;
      RECT 76.463 72.604 76.513 80.025 ;
      RECT 69.149 79.918 76.559 79.979 ;
      RECT 76.509 72.558 76.559 79.979 ;
      RECT 69.195 79.872 76.605 79.933 ;
      RECT 76.555 72.512 76.605 79.933 ;
      RECT 69.241 79.826 76.651 79.887 ;
      RECT 76.601 72.466 76.651 79.887 ;
      RECT 69.287 79.78 76.697 79.841 ;
      RECT 76.647 72.42 76.697 79.841 ;
      RECT 69.333 79.734 76.743 79.795 ;
      RECT 76.693 72.374 76.743 79.795 ;
      RECT 69.379 79.688 76.789 79.749 ;
      RECT 76.739 72.328 76.789 79.749 ;
      RECT 69.425 79.642 76.825 79.708 ;
      RECT 71.035 78.032 71.085 85.453 ;
      RECT 69.471 79.596 76.871 79.667 ;
      RECT 76.785 72.282 76.871 79.667 ;
      RECT 69.517 79.55 76.917 79.621 ;
      RECT 76.831 72.236 76.917 79.621 ;
      RECT 69.563 79.504 76.963 79.575 ;
      RECT 76.877 72.19 76.963 79.575 ;
      RECT 69.609 79.458 77.009 79.529 ;
      RECT 76.923 72.144 77.009 79.529 ;
      RECT 69.655 79.412 77.055 79.483 ;
      RECT 76.969 72.098 77.055 79.483 ;
      RECT 69.701 79.366 77.101 79.437 ;
      RECT 77.015 72.052 77.101 79.437 ;
      RECT 69.747 79.32 77.147 79.391 ;
      RECT 77.061 72.006 77.147 79.391 ;
      RECT 69.793 79.274 77.193 79.345 ;
      RECT 77.107 71.96 77.193 79.345 ;
      RECT 69.839 79.228 77.239 79.299 ;
      RECT 77.153 71.914 77.239 79.299 ;
      RECT 69.885 79.182 77.285 79.253 ;
      RECT 77.199 71.868 77.285 79.253 ;
      RECT 69.931 79.136 77.331 79.207 ;
      RECT 77.245 71.822 77.331 79.207 ;
      RECT 69.977 79.09 77.377 79.161 ;
      RECT 77.291 71.776 77.377 79.161 ;
      RECT 70.023 79.044 77.423 79.115 ;
      RECT 77.337 71.73 77.423 79.115 ;
      RECT 70.069 78.998 77.469 79.069 ;
      RECT 77.383 71.684 77.469 79.069 ;
      RECT 70.115 78.952 77.515 79.023 ;
      RECT 77.429 71.638 77.515 79.023 ;
      RECT 70.161 78.906 77.561 78.977 ;
      RECT 77.475 71.592 77.561 78.977 ;
      RECT 70.207 78.86 77.607 78.931 ;
      RECT 77.521 71.546 77.607 78.931 ;
      RECT 70.253 78.814 77.653 78.885 ;
      RECT 77.567 71.5 77.653 78.885 ;
      RECT 70.299 78.768 77.699 78.839 ;
      RECT 77.613 71.454 77.699 78.839 ;
      RECT 70.345 78.722 77.745 78.793 ;
      RECT 77.659 71.408 77.745 78.793 ;
      RECT 70.391 78.676 77.791 78.747 ;
      RECT 77.705 71.362 77.791 78.747 ;
      RECT 70.437 78.63 77.837 78.701 ;
      RECT 77.751 71.316 77.837 78.701 ;
      RECT 70.483 78.584 77.883 78.655 ;
      RECT 77.797 71.27 77.883 78.655 ;
      RECT 70.529 78.538 77.929 78.609 ;
      RECT 77.843 71.224 77.929 78.609 ;
      RECT 70.575 78.492 77.975 78.563 ;
      RECT 77.889 71.178 77.975 78.563 ;
      RECT 70.621 78.446 78.021 78.517 ;
      RECT 77.935 71.132 78.021 78.517 ;
      RECT 70.667 78.4 78.067 78.471 ;
      RECT 77.981 71.086 78.067 78.471 ;
      RECT 70.713 78.354 78.113 78.425 ;
      RECT 78.027 71.04 78.113 78.425 ;
      RECT 70.759 78.308 78.159 78.379 ;
      RECT 78.073 70.994 78.159 78.379 ;
      RECT 70.805 78.262 78.205 78.333 ;
      RECT 78.119 70.948 78.205 78.333 ;
      RECT 70.851 78.216 78.251 78.287 ;
      RECT 78.165 70.902 78.251 78.287 ;
      RECT 70.897 78.17 78.297 78.241 ;
      RECT 78.211 70.856 78.297 78.241 ;
      RECT 70.943 78.124 78.343 78.195 ;
      RECT 78.257 70.81 78.343 78.195 ;
      RECT 70.989 78.078 78.389 78.149 ;
      RECT 78.303 70.764 78.389 78.149 ;
      RECT 78.349 70.718 78.435 78.103 ;
      RECT 78.395 70.672 78.481 78.057 ;
      RECT 78.441 70.626 78.527 78.011 ;
      RECT 78.487 70.58 78.573 77.965 ;
      RECT 78.533 70.534 78.619 77.919 ;
      RECT 78.579 70.488 78.665 77.873 ;
      RECT 78.625 70.442 78.711 77.827 ;
      RECT 78.671 70.396 78.757 77.781 ;
      RECT 78.717 70.35 78.803 77.735 ;
      RECT 78.763 70.304 78.849 77.689 ;
      RECT 78.809 70.258 78.895 77.643 ;
      RECT 78.855 70.212 78.941 77.597 ;
      RECT 78.901 70.166 78.987 77.551 ;
      RECT 78.947 70.12 79.033 77.505 ;
      RECT 78.993 70.074 79.079 77.459 ;
      RECT 79.039 70.028 79.125 77.413 ;
      RECT 79.085 69.982 79.171 77.367 ;
      RECT 79.131 69.936 79.217 77.321 ;
      RECT 79.177 69.89 79.263 77.275 ;
      RECT 79.223 69.844 79.309 77.229 ;
      RECT 79.269 69.798 79.355 77.183 ;
      RECT 79.315 69.752 79.401 77.137 ;
      RECT 79.361 69.706 79.447 77.091 ;
      RECT 79.407 69.66 79.493 77.045 ;
      RECT 79.453 69.614 79.539 76.999 ;
      RECT 79.499 69.568 79.585 76.953 ;
      RECT 79.545 69.522 79.631 76.907 ;
      RECT 79.591 69.476 79.677 76.861 ;
      RECT 79.637 69.43 79.723 76.815 ;
      RECT 79.683 69.384 79.769 76.769 ;
      RECT 79.729 69.338 79.815 76.723 ;
      RECT 79.775 69.292 79.861 76.677 ;
      RECT 79.821 69.246 79.907 76.631 ;
      RECT 79.867 69.2 79.953 76.585 ;
      RECT 79.913 69.154 79.999 76.539 ;
      RECT 79.959 69.108 80.045 76.493 ;
      RECT 80.005 69.062 80.091 76.447 ;
      RECT 80.051 69.016 80.137 76.401 ;
      RECT 80.097 68.97 80.183 76.355 ;
      RECT 80.143 68.924 80.229 76.309 ;
      RECT 80.189 68.878 80.275 76.263 ;
      RECT 80.235 68.832 80.321 76.217 ;
      RECT 80.281 68.786 80.367 76.171 ;
      RECT 80.327 68.74 80.413 76.125 ;
      RECT 80.373 68.694 80.459 76.079 ;
      RECT 80.419 68.648 80.505 76.033 ;
      RECT 80.465 68.602 80.551 75.987 ;
      RECT 80.511 68.556 80.597 75.941 ;
      RECT 80.557 68.51 80.643 75.895 ;
      RECT 80.603 68.464 80.689 75.849 ;
      RECT 80.649 68.418 80.735 75.803 ;
      RECT 80.695 68.372 80.781 75.757 ;
      RECT 80.741 68.326 80.827 75.711 ;
      RECT 80.787 68.28 80.873 75.665 ;
      RECT 80.833 68.234 80.919 75.619 ;
      RECT 80.879 68.188 80.965 75.573 ;
      RECT 80.925 68.142 81.011 75.527 ;
      RECT 80.971 68.096 81.057 75.481 ;
      RECT 81.017 68.05 81.103 75.435 ;
      RECT 81.063 68.004 81.149 75.389 ;
      RECT 81.109 67.958 81.195 75.343 ;
      RECT 81.155 67.912 81.241 75.297 ;
      RECT 81.201 67.866 81.287 75.251 ;
      RECT 81.247 67.82 81.333 75.205 ;
      RECT 81.293 67.774 81.379 75.159 ;
      RECT 81.339 67.728 81.425 75.113 ;
      RECT 81.385 67.682 81.471 75.067 ;
      RECT 81.431 67.636 81.517 75.021 ;
      RECT 81.477 67.59 81.563 74.975 ;
      RECT 81.523 67.544 81.609 74.929 ;
      RECT 81.569 67.498 81.655 74.883 ;
      RECT 81.615 67.452 81.701 74.837 ;
      RECT 81.661 67.406 81.747 74.791 ;
      RECT 81.707 67.36 81.793 74.745 ;
      RECT 81.753 67.314 81.839 74.699 ;
      RECT 81.799 67.268 81.885 74.653 ;
      RECT 81.845 67.222 81.931 74.607 ;
      RECT 81.891 67.176 81.977 74.561 ;
      RECT 81.937 67.13 82.023 74.515 ;
      RECT 81.983 67.084 82.069 74.469 ;
      RECT 82.029 67.038 82.115 74.423 ;
      RECT 82.075 66.992 82.161 74.377 ;
      RECT 82.121 66.946 82.207 74.331 ;
      RECT 82.167 66.9 82.253 74.285 ;
      RECT 82.213 66.854 82.299 74.239 ;
      RECT 82.259 66.808 82.345 74.193 ;
      RECT 82.305 66.762 82.391 74.147 ;
      RECT 82.351 66.716 82.437 74.101 ;
      RECT 82.397 66.67 82.483 74.055 ;
      RECT 82.443 66.624 82.529 74.009 ;
      RECT 82.489 66.578 82.575 73.963 ;
      RECT 82.535 66.532 82.621 73.917 ;
      RECT 82.581 66.486 82.667 73.871 ;
      RECT 82.627 66.44 82.713 73.825 ;
      RECT 82.673 66.394 82.759 73.779 ;
      RECT 82.719 66.348 82.805 73.733 ;
      RECT 82.765 66.302 82.851 73.687 ;
      RECT 82.811 66.256 82.897 73.641 ;
      RECT 82.903 66.171 82.943 73.595 ;
      RECT 82.935 66.132 82.989 73.549 ;
      RECT 82.981 66.086 83.035 73.503 ;
      RECT 83.027 66.04 83.081 73.457 ;
      RECT 83.073 65.994 83.127 73.411 ;
      RECT 83.119 65.948 83.173 73.365 ;
      RECT 83.165 65.902 83.219 73.319 ;
      RECT 83.211 65.856 83.265 73.273 ;
      RECT 83.257 65.81 83.311 73.227 ;
      RECT 83.303 65.764 83.357 73.181 ;
      RECT 83.349 65.718 83.403 73.135 ;
      RECT 83.395 65.672 83.449 73.089 ;
      RECT 83.441 65.626 83.495 73.043 ;
      RECT 83.487 65.58 83.541 72.997 ;
      RECT 83.533 65.534 83.587 72.951 ;
      RECT 83.579 65.488 83.633 72.905 ;
      RECT 83.625 65.442 83.679 72.859 ;
      RECT 83.671 65.396 83.725 72.813 ;
      RECT 83.717 65.35 83.771 72.767 ;
      RECT 83.763 65.304 83.817 72.721 ;
      RECT 83.809 65.258 83.863 72.675 ;
      RECT 83.855 65.212 83.909 72.629 ;
      RECT 83.901 65.166 83.955 72.583 ;
      RECT 83.947 65.12 84.001 72.537 ;
      RECT 83.993 65.074 84.047 72.491 ;
      RECT 84.039 65.028 84.093 72.445 ;
      RECT 84.085 64.982 84.139 72.399 ;
      RECT 84.131 64.936 84.185 72.353 ;
      RECT 84.177 64.89 84.231 72.307 ;
      RECT 84.223 64.844 84.277 72.261 ;
      RECT 84.269 64.798 84.323 72.215 ;
      RECT 84.315 64.752 84.369 72.169 ;
      RECT 84.361 64.706 84.415 72.123 ;
      RECT 84.407 64.66 84.461 72.077 ;
      RECT 84.453 64.614 84.507 72.031 ;
      RECT 84.499 64.568 84.553 71.985 ;
      RECT 84.545 64.522 84.599 71.939 ;
      RECT 84.591 64.476 84.645 71.893 ;
      RECT 84.637 64.43 84.691 71.847 ;
      RECT 84.683 64.384 84.737 71.801 ;
      RECT 84.729 64.338 84.783 71.755 ;
      RECT 84.775 64.292 84.829 71.709 ;
      RECT 84.821 64.246 84.875 71.663 ;
      RECT 84.867 64.2 84.921 71.617 ;
      RECT 84.913 64.154 84.967 71.571 ;
      RECT 84.959 64.108 85.013 71.525 ;
      RECT 85.005 64.062 85.059 71.479 ;
      RECT 85.051 64.016 85.105 71.433 ;
      RECT 85.097 63.97 85.151 71.387 ;
      RECT 85.143 63.924 85.197 71.341 ;
      RECT 85.189 63.878 85.243 71.295 ;
      RECT 85.235 63.832 85.289 71.249 ;
      RECT 85.281 63.786 85.335 71.203 ;
      RECT 85.327 63.74 85.381 71.157 ;
      RECT 85.373 63.696 85.427 71.111 ;
      RECT 85.415 63.675 85.473 71.065 ;
      RECT 82.857 66.21 82.943 73.595 ;
      RECT 85.415 63.675 85.519 71.019 ;
      RECT 85.415 63.675 85.565 70.973 ;
      RECT 85.415 63.675 85.611 70.927 ;
      RECT 85.415 63.675 85.657 70.881 ;
      RECT 85.415 63.675 85.703 70.835 ;
      RECT 85.415 63.675 85.749 70.789 ;
      RECT 85.415 63.675 85.795 70.743 ;
      RECT 85.415 63.675 85.841 70.697 ;
      RECT 85.415 63.675 85.887 70.651 ;
      RECT 85.415 63.675 85.933 70.605 ;
      RECT 85.415 63.675 85.979 70.559 ;
      RECT 85.415 63.675 86.025 70.513 ;
      RECT 85.415 63.675 86.071 70.467 ;
      RECT 85.415 63.675 86.117 70.421 ;
      RECT 85.415 63.675 86.163 70.375 ;
      RECT 85.415 63.675 86.209 70.329 ;
      RECT 85.415 63.675 86.255 70.283 ;
      RECT 85.415 63.675 86.301 70.237 ;
      RECT 85.415 63.675 86.347 70.191 ;
      RECT 85.415 63.675 86.393 70.145 ;
      RECT 85.415 63.675 86.439 70.099 ;
      RECT 85.415 63.675 86.485 70.053 ;
      RECT 85.415 63.675 86.531 70.007 ;
      RECT 85.415 63.675 86.577 69.961 ;
      RECT 85.415 63.675 86.623 69.915 ;
      RECT 85.415 63.675 86.669 69.869 ;
      RECT 85.415 63.675 86.715 69.823 ;
      RECT 85.415 63.675 86.761 69.777 ;
      RECT 85.415 63.675 86.807 69.731 ;
      RECT 85.415 63.675 86.853 69.685 ;
      RECT 85.415 63.675 86.899 69.639 ;
      RECT 85.415 63.675 86.945 69.593 ;
      RECT 85.415 63.675 86.991 69.547 ;
      RECT 85.415 63.675 87.037 69.501 ;
      RECT 85.415 63.675 87.083 69.455 ;
      RECT 85.415 63.675 87.129 69.409 ;
      RECT 85.415 63.675 87.175 69.363 ;
      RECT 85.415 63.675 87.221 69.317 ;
      RECT 85.415 63.675 87.267 69.271 ;
      RECT 85.415 63.675 87.313 69.225 ;
      RECT 85.415 63.675 87.359 69.179 ;
      RECT 85.415 63.675 87.405 69.133 ;
      RECT 85.415 63.675 87.451 69.087 ;
      RECT 85.415 63.675 87.497 69.041 ;
      RECT 85.415 63.675 87.543 68.995 ;
      RECT 85.415 63.675 87.589 68.949 ;
      RECT 85.415 63.675 87.635 68.903 ;
      RECT 85.415 63.675 87.681 68.857 ;
      RECT 85.415 63.675 87.727 68.811 ;
      RECT 85.415 63.675 87.773 68.765 ;
      RECT 85.415 63.675 87.819 68.719 ;
      RECT 85.415 63.675 87.865 68.673 ;
      RECT 85.415 63.675 87.911 68.627 ;
      RECT 85.415 63.675 87.957 68.581 ;
      RECT 85.415 63.675 88.003 68.535 ;
      RECT 85.415 63.675 88.049 68.489 ;
      RECT 85.415 63.675 88.095 68.443 ;
      RECT 85.415 63.675 88.141 68.397 ;
      RECT 80.741 68.326 88.187 68.351 ;
      RECT 85.415 63.675 88.19 68.326 ;
      RECT 85.415 63.675 110 68.325 ;
      RECT 77.175 92.037 78.325 110 ;
      RECT 77.175 92.037 78.371 92.272 ;
      RECT 77.175 92.037 78.417 92.226 ;
      RECT 77.175 92.037 78.463 92.18 ;
      RECT 77.175 92.037 78.509 92.134 ;
      RECT 77.175 92.037 78.555 92.088 ;
      RECT 77.221 91.991 78.601 92.042 ;
      RECT 77.267 91.945 78.647 91.996 ;
      RECT 77.313 91.899 78.693 91.95 ;
      RECT 77.359 91.853 78.739 91.904 ;
      RECT 77.405 91.807 78.785 91.858 ;
      RECT 77.451 91.761 78.831 91.812 ;
      RECT 77.497 91.715 78.877 91.766 ;
      RECT 77.543 91.669 78.923 91.72 ;
      RECT 77.589 91.623 78.969 91.674 ;
      RECT 77.635 91.577 79.015 91.628 ;
      RECT 77.681 91.531 79.061 91.582 ;
      RECT 77.727 91.485 79.107 91.536 ;
      RECT 77.773 91.439 79.153 91.49 ;
      RECT 77.819 91.393 79.199 91.444 ;
      RECT 77.865 91.347 79.245 91.398 ;
      RECT 77.911 91.301 79.291 91.352 ;
      RECT 77.957 91.255 79.337 91.306 ;
      RECT 78.003 91.209 79.383 91.26 ;
      RECT 78.049 91.163 79.429 91.214 ;
      RECT 78.095 91.117 79.475 91.168 ;
      RECT 78.141 91.071 79.521 91.122 ;
      RECT 78.187 91.025 79.567 91.076 ;
      RECT 78.233 90.979 79.613 91.03 ;
      RECT 78.279 90.933 79.659 90.984 ;
      RECT 78.325 90.887 79.705 90.938 ;
      RECT 78.371 90.841 79.751 90.892 ;
      RECT 78.417 90.795 79.797 90.846 ;
      RECT 78.463 90.749 79.843 90.8 ;
      RECT 78.509 90.703 79.889 90.754 ;
      RECT 78.555 90.657 79.935 90.708 ;
      RECT 78.601 90.611 79.981 90.662 ;
      RECT 78.647 90.565 80.027 90.616 ;
      RECT 78.693 90.519 80.073 90.57 ;
      RECT 78.739 90.473 80.119 90.524 ;
      RECT 78.785 90.427 80.165 90.478 ;
      RECT 78.831 90.381 80.211 90.432 ;
      RECT 78.877 90.335 80.257 90.386 ;
      RECT 78.923 90.289 80.303 90.34 ;
      RECT 78.969 90.243 80.349 90.294 ;
      RECT 79.015 90.197 80.395 90.248 ;
      RECT 79.061 90.151 80.441 90.202 ;
      RECT 79.107 90.105 80.487 90.156 ;
      RECT 79.153 90.059 80.533 90.11 ;
      RECT 79.199 90.013 80.579 90.064 ;
      RECT 79.245 89.967 80.625 90.018 ;
      RECT 79.291 89.921 80.671 89.972 ;
      RECT 79.337 89.875 80.717 89.926 ;
      RECT 79.383 89.829 80.763 89.88 ;
      RECT 79.429 89.783 80.809 89.834 ;
      RECT 79.475 89.737 80.855 89.788 ;
      RECT 79.521 89.691 80.901 89.742 ;
      RECT 79.567 89.645 80.947 89.696 ;
      RECT 79.613 89.599 80.993 89.65 ;
      RECT 79.659 89.553 81.039 89.604 ;
      RECT 79.705 89.507 81.085 89.558 ;
      RECT 79.751 89.461 81.131 89.512 ;
      RECT 79.797 89.415 81.177 89.466 ;
      RECT 79.843 89.369 81.223 89.42 ;
      RECT 79.889 89.323 81.269 89.374 ;
      RECT 79.935 89.277 81.315 89.328 ;
      RECT 79.981 89.231 81.361 89.282 ;
      RECT 80.027 89.185 81.407 89.236 ;
      RECT 80.073 89.139 81.453 89.19 ;
      RECT 80.119 89.093 81.499 89.144 ;
      RECT 80.165 89.047 81.545 89.098 ;
      RECT 80.211 89.001 81.591 89.052 ;
      RECT 80.257 88.955 81.637 89.006 ;
      RECT 80.303 88.909 81.683 88.96 ;
      RECT 80.349 88.863 81.729 88.914 ;
      RECT 80.395 88.817 81.775 88.868 ;
      RECT 80.441 88.771 81.821 88.822 ;
      RECT 80.487 88.725 81.867 88.776 ;
      RECT 80.533 88.679 81.913 88.73 ;
      RECT 80.579 88.633 81.959 88.684 ;
      RECT 80.625 88.587 82.005 88.638 ;
      RECT 80.671 88.541 82.051 88.592 ;
      RECT 80.717 88.495 82.097 88.546 ;
      RECT 80.763 88.449 82.143 88.5 ;
      RECT 80.809 88.403 82.189 88.454 ;
      RECT 80.855 88.357 82.235 88.408 ;
      RECT 80.901 88.311 82.281 88.362 ;
      RECT 80.947 88.265 82.327 88.316 ;
      RECT 80.993 88.219 82.373 88.27 ;
      RECT 81.039 88.173 82.419 88.224 ;
      RECT 81.085 88.127 82.465 88.178 ;
      RECT 81.131 88.081 82.511 88.132 ;
      RECT 81.177 88.035 82.557 88.086 ;
      RECT 81.223 87.989 82.603 88.04 ;
      RECT 81.269 87.943 82.649 87.994 ;
      RECT 81.315 87.897 82.695 87.948 ;
      RECT 81.361 87.851 82.741 87.902 ;
      RECT 81.407 87.805 82.787 87.856 ;
      RECT 81.453 87.759 82.833 87.81 ;
      RECT 81.499 87.713 82.879 87.764 ;
      RECT 81.545 87.667 82.925 87.718 ;
      RECT 81.591 87.621 82.971 87.672 ;
      RECT 81.637 87.575 83.017 87.626 ;
      RECT 81.683 87.529 83.063 87.58 ;
      RECT 81.729 87.483 83.109 87.534 ;
      RECT 81.775 87.437 83.155 87.488 ;
      RECT 81.821 87.391 83.201 87.442 ;
      RECT 81.867 87.345 83.247 87.396 ;
      RECT 81.913 87.299 83.293 87.35 ;
      RECT 81.959 87.253 83.339 87.304 ;
      RECT 82.005 87.207 83.385 87.258 ;
      RECT 82.051 87.161 83.431 87.212 ;
      RECT 82.097 87.115 83.477 87.166 ;
      RECT 82.143 87.069 83.523 87.12 ;
      RECT 82.189 87.023 83.569 87.074 ;
      RECT 82.235 86.977 83.615 87.028 ;
      RECT 82.281 86.931 83.661 86.982 ;
      RECT 82.327 86.885 83.707 86.936 ;
      RECT 82.373 86.839 83.753 86.89 ;
      RECT 82.419 86.793 83.799 86.844 ;
      RECT 82.465 86.747 83.845 86.798 ;
      RECT 82.511 86.701 83.891 86.752 ;
      RECT 82.557 86.655 83.937 86.706 ;
      RECT 82.603 86.609 83.983 86.66 ;
      RECT 82.649 86.563 84.029 86.614 ;
      RECT 82.695 86.517 84.075 86.568 ;
      RECT 82.741 86.471 84.121 86.522 ;
      RECT 82.787 86.425 84.167 86.476 ;
      RECT 82.833 86.379 84.213 86.43 ;
      RECT 82.879 86.333 84.259 86.384 ;
      RECT 82.925 86.287 84.305 86.338 ;
      RECT 82.971 86.241 84.351 86.292 ;
      RECT 83.017 86.195 84.397 86.246 ;
      RECT 83.063 86.149 84.443 86.2 ;
      RECT 83.109 86.103 84.489 86.154 ;
      RECT 83.155 86.057 84.535 86.108 ;
      RECT 83.201 86.011 84.581 86.062 ;
      RECT 83.247 85.965 84.627 86.016 ;
      RECT 83.293 85.919 84.673 85.97 ;
      RECT 83.339 85.873 84.719 85.924 ;
      RECT 83.385 85.827 84.765 85.878 ;
      RECT 83.431 85.781 84.811 85.832 ;
      RECT 83.477 85.735 84.857 85.786 ;
      RECT 83.523 85.689 84.903 85.74 ;
      RECT 83.569 85.643 84.949 85.694 ;
      RECT 83.615 85.597 84.995 85.648 ;
      RECT 83.661 85.551 85.041 85.602 ;
      RECT 83.707 85.505 85.087 85.556 ;
      RECT 83.753 85.459 85.133 85.51 ;
      RECT 83.799 85.413 85.179 85.464 ;
      RECT 83.845 85.367 85.225 85.418 ;
      RECT 83.891 85.321 85.271 85.372 ;
      RECT 83.937 85.275 85.317 85.326 ;
      RECT 83.983 85.229 85.363 85.28 ;
      RECT 84.029 85.183 85.409 85.234 ;
      RECT 84.075 85.137 85.455 85.188 ;
      RECT 84.121 85.091 85.501 85.142 ;
      RECT 84.167 85.045 85.547 85.096 ;
      RECT 84.213 84.999 85.593 85.05 ;
      RECT 84.259 84.953 85.639 85.004 ;
      RECT 84.305 84.907 85.685 84.958 ;
      RECT 84.351 84.861 85.731 84.912 ;
      RECT 84.397 84.815 85.777 84.866 ;
      RECT 84.443 84.769 85.823 84.82 ;
      RECT 84.489 84.723 85.869 84.774 ;
      RECT 84.535 84.677 85.915 84.728 ;
      RECT 84.581 84.631 85.961 84.682 ;
      RECT 84.627 84.585 86.007 84.636 ;
      RECT 84.673 84.539 86.053 84.59 ;
      RECT 84.719 84.493 86.099 84.544 ;
      RECT 84.765 84.447 86.145 84.498 ;
      RECT 84.811 84.401 86.191 84.452 ;
      RECT 84.857 84.355 86.237 84.406 ;
      RECT 84.903 84.309 86.283 84.36 ;
      RECT 84.949 84.263 86.329 84.314 ;
      RECT 84.995 84.217 86.375 84.268 ;
      RECT 85.041 84.171 86.421 84.222 ;
      RECT 85.087 84.125 86.467 84.176 ;
      RECT 85.133 84.079 86.513 84.13 ;
      RECT 85.179 84.033 86.559 84.084 ;
      RECT 85.225 83.987 86.605 84.038 ;
      RECT 85.271 83.941 86.651 83.992 ;
      RECT 85.317 83.895 86.697 83.946 ;
      RECT 85.363 83.849 86.743 83.9 ;
      RECT 85.409 83.803 86.789 83.854 ;
      RECT 85.455 83.757 86.835 83.808 ;
      RECT 85.501 83.711 86.881 83.762 ;
      RECT 85.547 83.665 86.927 83.716 ;
      RECT 85.593 83.619 86.973 83.67 ;
      RECT 85.639 83.573 87.019 83.624 ;
      RECT 85.685 83.527 87.065 83.578 ;
      RECT 85.731 83.481 87.111 83.532 ;
      RECT 85.777 83.435 87.157 83.486 ;
      RECT 85.823 83.389 87.203 83.44 ;
      RECT 85.869 83.343 87.249 83.394 ;
      RECT 85.915 83.297 87.295 83.348 ;
      RECT 85.961 83.251 87.341 83.302 ;
      RECT 86.007 83.205 87.387 83.256 ;
      RECT 86.053 83.159 87.433 83.21 ;
      RECT 86.099 83.113 87.479 83.164 ;
      RECT 86.145 83.067 87.525 83.118 ;
      RECT 86.191 83.021 87.571 83.072 ;
      RECT 86.237 82.975 87.617 83.026 ;
      RECT 86.283 82.929 87.663 82.98 ;
      RECT 86.329 82.883 87.709 82.934 ;
      RECT 86.375 82.837 87.755 82.888 ;
      RECT 86.421 82.791 87.801 82.842 ;
      RECT 86.467 82.745 87.847 82.796 ;
      RECT 86.513 82.699 87.893 82.75 ;
      RECT 86.559 82.653 87.939 82.704 ;
      RECT 86.605 82.607 87.985 82.658 ;
      RECT 86.651 82.561 88.031 82.612 ;
      RECT 86.697 82.515 88.077 82.566 ;
      RECT 86.743 82.469 88.123 82.52 ;
      RECT 86.789 82.423 88.169 82.474 ;
      RECT 86.835 82.377 88.215 82.428 ;
      RECT 86.881 82.331 88.261 82.382 ;
      RECT 86.927 82.285 88.307 82.336 ;
      RECT 86.973 82.239 88.353 82.29 ;
      RECT 87.019 82.193 88.399 82.244 ;
      RECT 87.065 82.147 88.445 82.198 ;
      RECT 87.111 82.101 88.491 82.152 ;
      RECT 87.157 82.055 88.537 82.106 ;
      RECT 87.203 82.009 88.583 82.06 ;
      RECT 88.537 80.697 88.583 82.06 ;
      RECT 87.249 81.963 88.629 82.014 ;
      RECT 87.295 81.917 88.675 81.968 ;
      RECT 87.341 81.871 88.721 81.922 ;
      RECT 87.387 81.825 88.767 81.876 ;
      RECT 87.433 81.779 88.813 81.83 ;
      RECT 87.479 81.733 88.859 81.784 ;
      RECT 87.525 81.687 88.905 81.738 ;
      RECT 87.571 81.641 88.951 81.692 ;
      RECT 87.617 81.595 88.997 81.646 ;
      RECT 87.663 81.549 89.043 81.6 ;
      RECT 87.709 81.503 89.089 81.554 ;
      RECT 87.755 81.457 89.135 81.508 ;
      RECT 87.801 81.411 89.181 81.462 ;
      RECT 87.847 81.365 89.227 81.416 ;
      RECT 87.893 81.319 89.273 81.37 ;
      RECT 87.939 81.273 89.319 81.324 ;
      RECT 87.939 81.273 89.325 81.298 ;
      RECT 87.985 81.227 89.371 81.272 ;
      RECT 88.031 81.181 89.417 81.226 ;
      RECT 88.077 81.135 89.463 81.18 ;
      RECT 88.123 81.089 89.509 81.134 ;
      RECT 88.169 81.043 89.555 81.088 ;
      RECT 88.215 80.997 89.601 81.042 ;
      RECT 88.261 80.951 89.647 80.996 ;
      RECT 88.307 80.905 89.693 80.95 ;
      RECT 88.353 80.859 89.739 80.904 ;
      RECT 88.399 80.813 89.785 80.858 ;
      RECT 88.445 80.767 89.831 80.812 ;
      RECT 88.491 80.721 89.877 80.766 ;
      RECT 88.54 80.672 89.923 80.72 ;
      RECT 89.874 79.338 89.923 80.72 ;
      RECT 88.586 80.626 89.969 80.674 ;
      RECT 89.92 79.292 89.969 80.674 ;
      RECT 88.632 80.58 90.015 80.628 ;
      RECT 89.966 79.246 90.015 80.628 ;
      RECT 88.678 80.534 90.061 80.582 ;
      RECT 90.012 79.2 90.061 80.582 ;
      RECT 88.724 80.488 90.107 80.536 ;
      RECT 90.058 79.154 90.107 80.536 ;
      RECT 88.77 80.442 90.153 80.49 ;
      RECT 90.104 79.108 90.153 80.49 ;
      RECT 88.816 80.396 90.199 80.444 ;
      RECT 90.15 79.062 90.199 80.444 ;
      RECT 88.862 80.35 90.245 80.398 ;
      RECT 90.196 79.016 90.245 80.398 ;
      RECT 88.908 80.304 90.291 80.352 ;
      RECT 90.242 78.97 90.291 80.352 ;
      RECT 88.954 80.258 90.337 80.306 ;
      RECT 90.288 78.924 90.337 80.306 ;
      RECT 89 80.212 90.383 80.26 ;
      RECT 90.334 78.878 90.383 80.26 ;
      RECT 89.046 80.166 90.429 80.214 ;
      RECT 90.38 78.832 90.429 80.214 ;
      RECT 89.092 80.12 90.475 80.168 ;
      RECT 90.426 78.786 90.475 80.168 ;
      RECT 89.138 80.074 90.521 80.122 ;
      RECT 90.472 78.74 90.521 80.122 ;
      RECT 89.184 80.028 90.567 80.076 ;
      RECT 90.518 78.694 90.567 80.076 ;
      RECT 89.23 79.982 90.613 80.03 ;
      RECT 90.564 78.648 90.613 80.03 ;
      RECT 89.276 79.936 90.659 79.984 ;
      RECT 90.61 78.602 90.659 79.984 ;
      RECT 89.322 79.89 90.705 79.938 ;
      RECT 90.656 78.556 90.705 79.938 ;
      RECT 89.368 79.844 90.751 79.892 ;
      RECT 90.702 78.51 90.751 79.892 ;
      RECT 89.414 79.798 90.797 79.846 ;
      RECT 90.748 78.464 90.797 79.846 ;
      RECT 89.46 79.752 90.843 79.8 ;
      RECT 90.794 78.418 90.843 79.8 ;
      RECT 89.506 79.706 90.889 79.754 ;
      RECT 90.84 78.372 90.889 79.754 ;
      RECT 89.552 79.66 90.935 79.708 ;
      RECT 90.886 78.326 90.935 79.708 ;
      RECT 89.598 79.614 90.981 79.662 ;
      RECT 90.932 78.28 90.981 79.662 ;
      RECT 89.644 79.568 91.027 79.616 ;
      RECT 90.978 78.234 91.027 79.616 ;
      RECT 89.69 79.522 91.073 79.57 ;
      RECT 91.024 78.188 91.073 79.57 ;
      RECT 89.736 79.476 91.119 79.524 ;
      RECT 91.07 78.142 91.119 79.524 ;
      RECT 89.782 79.43 91.165 79.478 ;
      RECT 91.116 78.096 91.165 79.478 ;
      RECT 89.828 79.384 91.211 79.432 ;
      RECT 91.162 78.05 91.211 79.432 ;
      RECT 91.208 78.004 91.257 79.386 ;
      RECT 91.254 77.958 91.303 79.34 ;
      RECT 91.3 77.912 91.349 79.294 ;
      RECT 91.346 77.866 91.395 79.248 ;
      RECT 91.392 77.82 91.441 79.202 ;
      RECT 91.438 77.774 91.487 79.156 ;
      RECT 91.484 77.728 91.533 79.11 ;
      RECT 91.53 77.682 91.579 79.064 ;
      RECT 91.576 77.636 91.625 79.018 ;
      RECT 91.622 77.59 91.671 78.972 ;
      RECT 91.668 77.544 91.717 78.926 ;
      RECT 91.714 77.498 91.763 78.88 ;
      RECT 91.76 77.452 91.809 78.834 ;
      RECT 91.806 77.406 91.855 78.788 ;
      RECT 91.852 77.36 91.901 78.742 ;
      RECT 91.898 77.314 91.947 78.696 ;
      RECT 91.944 77.268 91.993 78.65 ;
      RECT 91.99 77.222 92.039 78.604 ;
      RECT 92.036 77.187 92.085 78.558 ;
      RECT 92.06 77.175 92.131 78.512 ;
      RECT 92.06 77.175 92.177 78.466 ;
      RECT 92.06 77.175 92.223 78.42 ;
      RECT 92.06 77.175 92.269 78.374 ;
      RECT 90.886 78.326 92.295 78.338 ;
      RECT 92.06 77.175 110 78.325 ;
      RECT 89.675 97.182 90.825 110 ;
      RECT 89.675 97.182 90.871 99.352 ;
      RECT 89.675 97.182 90.917 99.306 ;
      RECT 89.675 97.182 90.963 99.26 ;
      RECT 89.675 97.182 91.009 99.214 ;
      RECT 89.675 97.182 91.055 99.168 ;
      RECT 89.675 97.182 91.101 99.122 ;
      RECT 89.675 97.182 91.147 99.076 ;
      RECT 89.675 97.182 91.193 99.03 ;
      RECT 89.675 97.182 91.239 98.984 ;
      RECT 89.675 97.182 91.285 98.938 ;
      RECT 89.675 97.182 91.331 98.892 ;
      RECT 89.675 97.182 91.377 98.846 ;
      RECT 89.675 97.182 91.423 98.8 ;
      RECT 89.675 97.182 91.469 98.754 ;
      RECT 89.675 97.182 91.515 98.708 ;
      RECT 89.675 97.182 91.561 98.662 ;
      RECT 89.675 97.182 91.607 98.616 ;
      RECT 89.675 97.182 91.653 98.57 ;
      RECT 89.675 97.182 91.699 98.524 ;
      RECT 89.675 97.182 91.745 98.478 ;
      RECT 89.675 97.182 91.791 98.432 ;
      RECT 89.675 97.182 91.837 98.386 ;
      RECT 89.675 97.182 91.883 98.34 ;
      RECT 89.675 97.182 91.929 98.294 ;
      RECT 89.675 97.182 91.975 98.248 ;
      RECT 89.675 97.182 92.021 98.202 ;
      RECT 89.675 97.182 92.067 98.156 ;
      RECT 89.675 97.182 92.113 98.11 ;
      RECT 89.675 97.182 92.159 98.064 ;
      RECT 89.675 97.182 92.205 98.018 ;
      RECT 89.675 97.182 92.251 97.972 ;
      RECT 89.675 97.182 92.297 97.926 ;
      RECT 89.675 97.182 92.343 97.88 ;
      RECT 89.675 97.182 92.389 97.834 ;
      RECT 89.675 97.182 92.435 97.788 ;
      RECT 89.675 97.182 92.481 97.742 ;
      RECT 89.675 97.182 92.527 97.696 ;
      RECT 89.675 97.182 92.573 97.65 ;
      RECT 89.675 97.182 92.619 97.604 ;
      RECT 89.675 97.182 92.665 97.558 ;
      RECT 89.675 97.182 92.711 97.512 ;
      RECT 89.675 97.182 92.757 97.466 ;
      RECT 89.675 97.182 92.803 97.42 ;
      RECT 89.675 97.182 92.849 97.374 ;
      RECT 89.675 97.182 92.895 97.328 ;
      RECT 89.675 97.182 92.941 97.282 ;
      RECT 89.721 97.136 93.033 97.19 ;
      RECT 92.967 93.89 93.033 97.19 ;
      RECT 89.767 97.09 93.079 97.144 ;
      RECT 93.013 93.844 93.079 97.144 ;
      RECT 89.813 97.044 93.125 97.098 ;
      RECT 93.059 93.798 93.125 97.098 ;
      RECT 89.859 96.998 93.171 97.052 ;
      RECT 93.105 93.752 93.171 97.052 ;
      RECT 89.905 96.952 93.217 97.006 ;
      RECT 93.151 93.706 93.217 97.006 ;
      RECT 89.951 96.906 93.263 96.96 ;
      RECT 93.197 93.66 93.263 96.96 ;
      RECT 89.997 96.86 93.309 96.914 ;
      RECT 93.243 93.614 93.309 96.914 ;
      RECT 90.043 96.814 93.355 96.868 ;
      RECT 93.289 93.568 93.355 96.868 ;
      RECT 90.089 96.768 93.401 96.822 ;
      RECT 93.335 93.522 93.401 96.822 ;
      RECT 90.135 96.722 93.447 96.776 ;
      RECT 93.381 93.476 93.447 96.776 ;
      RECT 90.181 96.676 93.493 96.73 ;
      RECT 93.427 93.43 93.493 96.73 ;
      RECT 90.227 96.63 93.539 96.684 ;
      RECT 93.473 93.384 93.539 96.684 ;
      RECT 90.273 96.584 93.585 96.638 ;
      RECT 93.519 93.338 93.585 96.638 ;
      RECT 90.319 96.538 93.631 96.592 ;
      RECT 93.565 93.292 93.631 96.592 ;
      RECT 90.365 96.492 93.677 96.546 ;
      RECT 93.611 93.246 93.677 96.546 ;
      RECT 90.411 96.446 93.723 96.5 ;
      RECT 93.657 93.2 93.723 96.5 ;
      RECT 90.457 96.4 93.769 96.454 ;
      RECT 93.703 93.154 93.769 96.454 ;
      RECT 90.503 96.354 93.815 96.408 ;
      RECT 93.749 93.108 93.815 96.408 ;
      RECT 90.549 96.308 93.861 96.362 ;
      RECT 93.795 93.062 93.861 96.362 ;
      RECT 90.595 96.262 93.907 96.316 ;
      RECT 93.841 93.016 93.907 96.316 ;
      RECT 90.641 96.216 93.953 96.27 ;
      RECT 93.887 92.97 93.953 96.27 ;
      RECT 90.687 96.17 93.999 96.224 ;
      RECT 93.933 92.924 93.999 96.224 ;
      RECT 90.733 96.124 94.045 96.178 ;
      RECT 93.979 92.878 94.045 96.178 ;
      RECT 90.779 96.078 94.091 96.132 ;
      RECT 94.025 92.832 94.091 96.132 ;
      RECT 90.825 96.032 94.137 96.086 ;
      RECT 94.071 92.786 94.137 96.086 ;
      RECT 90.871 95.986 94.183 96.04 ;
      RECT 94.117 92.74 94.183 96.04 ;
      RECT 90.917 95.94 94.229 95.994 ;
      RECT 94.163 92.694 94.229 95.994 ;
      RECT 90.963 95.894 94.275 95.948 ;
      RECT 94.209 92.648 94.275 95.948 ;
      RECT 91.009 95.848 94.321 95.902 ;
      RECT 94.255 92.602 94.321 95.902 ;
      RECT 91.055 95.802 94.367 95.856 ;
      RECT 94.301 92.556 94.367 95.856 ;
      RECT 91.101 95.756 94.413 95.81 ;
      RECT 94.347 92.51 94.413 95.81 ;
      RECT 91.147 95.71 94.459 95.764 ;
      RECT 94.393 92.464 94.459 95.764 ;
      RECT 91.193 95.664 94.505 95.718 ;
      RECT 94.439 92.418 94.505 95.718 ;
      RECT 91.239 95.618 94.551 95.672 ;
      RECT 94.485 92.372 94.551 95.672 ;
      RECT 91.285 95.572 94.597 95.626 ;
      RECT 94.531 92.326 94.597 95.626 ;
      RECT 91.331 95.526 94.643 95.58 ;
      RECT 94.577 92.28 94.643 95.58 ;
      RECT 91.377 95.48 94.689 95.534 ;
      RECT 94.623 92.234 94.689 95.534 ;
      RECT 91.423 95.434 94.735 95.488 ;
      RECT 94.669 92.188 94.735 95.488 ;
      RECT 91.469 95.388 94.781 95.442 ;
      RECT 94.715 92.142 94.781 95.442 ;
      RECT 91.515 95.342 94.827 95.396 ;
      RECT 94.761 92.096 94.827 95.396 ;
      RECT 91.561 95.296 94.873 95.35 ;
      RECT 94.807 92.05 94.873 95.35 ;
      RECT 91.607 95.25 94.919 95.304 ;
      RECT 94.853 92.004 94.919 95.304 ;
      RECT 91.653 95.204 94.965 95.258 ;
      RECT 94.899 91.958 94.965 95.258 ;
      RECT 91.699 95.158 95.011 95.212 ;
      RECT 94.945 91.912 95.011 95.212 ;
      RECT 91.745 95.112 95.057 95.166 ;
      RECT 94.991 91.866 95.057 95.166 ;
      RECT 91.791 95.066 95.103 95.12 ;
      RECT 95.037 91.82 95.103 95.12 ;
      RECT 91.837 95.02 95.149 95.074 ;
      RECT 95.083 91.774 95.149 95.074 ;
      RECT 91.883 94.974 95.195 95.028 ;
      RECT 95.129 91.728 95.195 95.028 ;
      RECT 91.929 94.928 95.241 94.982 ;
      RECT 95.175 91.682 95.241 94.982 ;
      RECT 91.975 94.882 95.287 94.936 ;
      RECT 95.221 91.636 95.287 94.936 ;
      RECT 92.021 94.836 95.333 94.89 ;
      RECT 95.267 91.59 95.333 94.89 ;
      RECT 92.067 94.79 95.379 94.844 ;
      RECT 95.313 91.544 95.379 94.844 ;
      RECT 92.113 94.744 95.425 94.798 ;
      RECT 95.359 91.498 95.425 94.798 ;
      RECT 92.159 94.698 95.471 94.752 ;
      RECT 95.405 91.452 95.471 94.752 ;
      RECT 92.205 94.652 95.517 94.706 ;
      RECT 95.451 91.406 95.517 94.706 ;
      RECT 92.251 94.606 95.563 94.66 ;
      RECT 95.497 91.36 95.563 94.66 ;
      RECT 92.297 94.56 95.609 94.614 ;
      RECT 95.543 91.314 95.609 94.614 ;
      RECT 92.343 94.514 95.655 94.568 ;
      RECT 95.589 91.268 95.655 94.568 ;
      RECT 92.389 94.468 95.701 94.522 ;
      RECT 95.635 91.222 95.701 94.522 ;
      RECT 92.435 94.422 95.747 94.476 ;
      RECT 95.681 91.176 95.747 94.476 ;
      RECT 92.481 94.376 95.793 94.43 ;
      RECT 95.727 91.13 95.793 94.43 ;
      RECT 92.527 94.33 95.839 94.384 ;
      RECT 95.773 91.084 95.839 94.384 ;
      RECT 92.573 94.284 95.885 94.338 ;
      RECT 95.819 91.038 95.885 94.338 ;
      RECT 92.619 94.248 95.931 94.292 ;
      RECT 95.865 90.992 95.931 94.292 ;
      RECT 92.645 94.212 95.931 94.292 ;
      RECT 92.921 93.936 92.987 97.236 ;
      RECT 92.691 94.166 95.977 94.246 ;
      RECT 95.911 90.946 95.977 94.246 ;
      RECT 92.737 94.12 96.023 94.2 ;
      RECT 95.957 90.9 96.023 94.2 ;
      RECT 92.783 94.074 96.069 94.154 ;
      RECT 96.003 90.854 96.069 94.154 ;
      RECT 92.829 94.028 96.115 94.108 ;
      RECT 96.049 90.808 96.115 94.108 ;
      RECT 92.875 93.982 96.161 94.062 ;
      RECT 96.095 90.762 96.161 94.062 ;
      RECT 96.141 90.716 96.207 94.016 ;
      RECT 96.187 90.67 96.253 93.97 ;
      RECT 96.233 90.624 96.299 93.924 ;
      RECT 96.279 90.578 96.345 93.878 ;
      RECT 96.325 90.532 96.391 93.832 ;
      RECT 96.371 90.486 96.437 93.786 ;
      RECT 96.417 90.44 96.483 93.74 ;
      RECT 96.463 90.394 96.529 93.694 ;
      RECT 96.509 90.348 96.575 93.648 ;
      RECT 96.555 90.302 96.621 93.602 ;
      RECT 96.601 90.256 96.667 93.556 ;
      RECT 96.647 90.21 96.713 93.51 ;
      RECT 96.693 90.164 96.759 93.464 ;
      RECT 96.739 90.118 96.805 93.418 ;
      RECT 96.785 90.072 96.851 93.372 ;
      RECT 96.831 90.026 96.897 93.326 ;
      RECT 96.877 89.98 96.943 93.28 ;
      RECT 96.923 89.934 96.989 93.234 ;
      RECT 96.969 89.888 97.035 93.188 ;
      RECT 97.015 89.842 97.081 93.142 ;
      RECT 97.061 89.796 97.127 93.096 ;
      RECT 97.107 89.75 97.173 93.05 ;
      RECT 97.199 89.678 97.219 93.004 ;
      RECT 97.205 89.675 97.265 92.958 ;
      RECT 97.153 89.704 97.219 93.004 ;
      RECT 97.205 89.675 97.311 92.912 ;
      RECT 97.205 89.675 97.357 92.866 ;
      RECT 97.205 89.675 97.403 92.82 ;
      RECT 97.205 89.675 97.449 92.774 ;
      RECT 97.205 89.675 97.495 92.728 ;
      RECT 97.205 89.675 97.541 92.682 ;
      RECT 97.205 89.675 97.587 92.636 ;
      RECT 97.205 89.675 97.633 92.59 ;
      RECT 97.205 89.675 97.679 92.544 ;
      RECT 97.205 89.675 97.725 92.498 ;
      RECT 97.205 89.675 97.771 92.452 ;
      RECT 94.485 92.372 97.817 92.406 ;
      RECT 97.205 89.675 97.825 92.379 ;
      RECT 97.205 89.675 97.871 92.352 ;
      RECT 97.205 89.675 97.917 92.306 ;
      RECT 97.205 89.675 97.963 92.26 ;
      RECT 97.205 89.675 98.009 92.214 ;
      RECT 97.205 89.675 98.055 92.168 ;
      RECT 97.205 89.675 98.101 92.122 ;
      RECT 97.205 89.675 98.147 92.076 ;
      RECT 97.205 89.675 98.193 92.03 ;
      RECT 97.205 89.675 98.239 91.984 ;
      RECT 97.205 89.675 98.285 91.938 ;
      RECT 97.205 89.675 98.331 91.892 ;
      RECT 97.205 89.675 98.377 91.846 ;
      RECT 97.205 89.675 98.423 91.8 ;
      RECT 97.205 89.675 98.469 91.754 ;
      RECT 97.205 89.675 98.515 91.708 ;
      RECT 97.205 89.675 98.561 91.662 ;
      RECT 97.205 89.675 98.607 91.616 ;
      RECT 97.205 89.675 98.653 91.57 ;
      RECT 97.205 89.675 98.699 91.524 ;
      RECT 97.205 89.675 98.745 91.478 ;
      RECT 97.205 89.675 98.791 91.432 ;
      RECT 97.205 89.675 98.837 91.386 ;
      RECT 97.205 89.675 98.883 91.34 ;
      RECT 97.205 89.675 98.929 91.294 ;
      RECT 97.205 89.675 98.975 91.248 ;
      RECT 97.205 89.675 99.021 91.202 ;
      RECT 97.205 89.675 99.067 91.156 ;
      RECT 97.205 89.675 99.113 91.11 ;
      RECT 97.205 89.675 99.159 91.064 ;
      RECT 97.205 89.675 99.205 91.018 ;
      RECT 97.205 89.675 99.251 90.972 ;
      RECT 97.205 89.675 99.297 90.926 ;
      RECT 97.205 89.675 99.343 90.88 ;
      RECT 96.049 90.808 99.375 90.841 ;
      RECT 97.205 89.675 110 90.825 ;
      RECT 98.175 102.602 99.325 110 ;
      RECT 98.175 102.602 99.371 103.642 ;
      RECT 98.175 102.602 99.417 103.596 ;
      RECT 98.175 102.602 99.463 103.55 ;
      RECT 98.175 102.602 99.509 103.504 ;
      RECT 98.175 102.602 99.555 103.458 ;
      RECT 98.175 102.602 99.601 103.412 ;
      RECT 98.175 102.602 99.647 103.366 ;
      RECT 98.175 102.602 99.693 103.32 ;
      RECT 98.175 102.602 99.739 103.274 ;
      RECT 98.175 102.602 99.785 103.228 ;
      RECT 98.175 102.602 99.831 103.182 ;
      RECT 98.175 102.602 99.877 103.136 ;
      RECT 98.175 102.602 99.923 103.09 ;
      RECT 98.175 102.602 99.969 103.044 ;
      RECT 98.175 102.602 100.015 102.998 ;
      RECT 98.175 102.602 100.061 102.952 ;
      RECT 98.175 102.602 100.107 102.906 ;
      RECT 98.175 102.602 100.153 102.86 ;
      RECT 98.175 102.602 100.199 102.814 ;
      RECT 98.175 102.602 100.245 102.768 ;
      RECT 98.175 102.602 100.291 102.722 ;
      RECT 98.175 102.602 100.337 102.676 ;
      RECT 98.221 102.556 100.383 102.63 ;
      RECT 100.323 100.454 100.383 102.63 ;
      RECT 98.267 102.51 100.429 102.584 ;
      RECT 100.369 100.408 100.429 102.584 ;
      RECT 98.313 102.464 100.475 102.538 ;
      RECT 100.415 100.362 100.475 102.538 ;
      RECT 98.359 102.418 100.521 102.492 ;
      RECT 100.461 100.316 100.521 102.492 ;
      RECT 98.405 102.372 100.567 102.446 ;
      RECT 100.507 100.27 100.567 102.446 ;
      RECT 98.451 102.326 100.613 102.4 ;
      RECT 100.553 100.224 100.613 102.4 ;
      RECT 98.497 102.28 100.659 102.354 ;
      RECT 100.599 100.178 100.659 102.354 ;
      RECT 98.543 102.234 100.705 102.308 ;
      RECT 100.645 100.132 100.705 102.308 ;
      RECT 98.589 102.188 100.751 102.262 ;
      RECT 100.691 100.086 100.751 102.262 ;
      RECT 98.635 102.142 100.797 102.216 ;
      RECT 100.737 100.04 100.797 102.216 ;
      RECT 98.681 102.096 100.843 102.17 ;
      RECT 100.783 99.994 100.843 102.17 ;
      RECT 98.727 102.05 100.889 102.124 ;
      RECT 100.829 99.948 100.889 102.124 ;
      RECT 98.773 102.004 100.935 102.078 ;
      RECT 100.875 99.902 100.935 102.078 ;
      RECT 98.819 101.958 100.981 102.032 ;
      RECT 100.921 99.856 100.981 102.032 ;
      RECT 98.865 101.912 101.027 101.986 ;
      RECT 100.967 99.81 101.027 101.986 ;
      RECT 98.911 101.866 101.073 101.94 ;
      RECT 101.013 99.764 101.073 101.94 ;
      RECT 98.957 101.82 101.119 101.894 ;
      RECT 101.059 99.718 101.119 101.894 ;
      RECT 99.003 101.774 101.165 101.848 ;
      RECT 101.105 99.672 101.165 101.848 ;
      RECT 99.049 101.728 101.211 101.802 ;
      RECT 101.151 99.626 101.211 101.802 ;
      RECT 99.095 101.682 101.257 101.756 ;
      RECT 101.197 99.58 101.257 101.756 ;
      RECT 99.141 101.636 101.303 101.71 ;
      RECT 101.243 99.534 101.303 101.71 ;
      RECT 99.187 101.59 101.349 101.664 ;
      RECT 101.289 99.488 101.349 101.664 ;
      RECT 99.233 101.544 101.395 101.618 ;
      RECT 101.335 99.442 101.395 101.618 ;
      RECT 99.279 101.498 101.441 101.572 ;
      RECT 101.381 99.396 101.441 101.572 ;
      RECT 99.325 101.452 101.487 101.526 ;
      RECT 101.427 99.35 101.487 101.526 ;
      RECT 99.371 101.406 101.533 101.48 ;
      RECT 101.473 99.304 101.533 101.48 ;
      RECT 99.417 101.36 101.579 101.434 ;
      RECT 101.519 99.258 101.579 101.434 ;
      RECT 99.463 101.314 101.625 101.388 ;
      RECT 101.565 99.212 101.625 101.388 ;
      RECT 99.509 101.268 101.671 101.342 ;
      RECT 101.611 99.166 101.671 101.342 ;
      RECT 99.555 101.222 101.717 101.296 ;
      RECT 101.657 99.12 101.717 101.296 ;
      RECT 99.601 101.176 101.763 101.25 ;
      RECT 101.703 99.074 101.763 101.25 ;
      RECT 99.647 101.13 101.809 101.204 ;
      RECT 101.749 99.028 101.809 101.204 ;
      RECT 99.693 101.091 101.855 101.158 ;
      RECT 101.795 98.982 101.855 101.158 ;
      RECT 99.725 101.052 101.901 101.112 ;
      RECT 101.841 98.936 101.901 101.112 ;
      RECT 99.771 101.006 101.947 101.066 ;
      RECT 101.887 98.89 101.947 101.066 ;
      RECT 99.817 100.96 101.993 101.02 ;
      RECT 101.933 98.844 101.993 101.02 ;
      RECT 99.863 100.914 102.039 100.974 ;
      RECT 101.979 98.798 102.039 100.974 ;
      RECT 99.909 100.868 102.085 100.928 ;
      RECT 102.025 98.752 102.085 100.928 ;
      RECT 99.955 100.822 102.131 100.882 ;
      RECT 102.071 98.706 102.131 100.882 ;
      RECT 100.001 100.776 102.177 100.836 ;
      RECT 102.117 98.66 102.177 100.836 ;
      RECT 100.047 100.73 102.223 100.79 ;
      RECT 102.163 98.614 102.223 100.79 ;
      RECT 100.093 100.684 102.269 100.744 ;
      RECT 102.209 98.568 102.269 100.744 ;
      RECT 100.139 100.638 102.315 100.698 ;
      RECT 102.255 98.522 102.315 100.698 ;
      RECT 100.185 100.592 102.361 100.652 ;
      RECT 102.301 98.476 102.361 100.652 ;
      RECT 100.231 100.546 102.407 100.606 ;
      RECT 102.347 98.43 102.407 100.606 ;
      RECT 100.277 100.5 102.453 100.56 ;
      RECT 102.393 98.384 102.453 100.56 ;
      RECT 102.439 98.338 102.499 100.514 ;
      RECT 102.485 98.292 102.545 100.468 ;
      RECT 102.531 98.246 102.591 100.422 ;
      RECT 102.577 98.199 102.637 100.376 ;
      RECT 102.623 98.175 102.683 100.33 ;
      RECT 102.623 98.175 102.729 100.284 ;
      RECT 102.623 98.175 102.775 100.238 ;
      RECT 102.623 98.175 102.821 100.192 ;
      RECT 102.623 98.175 102.867 100.146 ;
      RECT 102.623 98.175 102.913 100.1 ;
      RECT 102.623 98.175 102.959 100.054 ;
      RECT 102.623 98.175 103.005 100.008 ;
      RECT 102.623 98.175 103.051 99.962 ;
      RECT 102.623 98.175 103.097 99.916 ;
      RECT 102.623 98.175 103.143 99.87 ;
      RECT 102.623 98.175 103.189 99.824 ;
      RECT 102.623 98.175 103.235 99.778 ;
      RECT 102.623 98.175 103.281 99.732 ;
      RECT 102.623 98.175 103.327 99.686 ;
      RECT 102.623 98.175 103.373 99.64 ;
      RECT 102.623 98.175 103.419 99.594 ;
      RECT 102.623 98.175 103.465 99.548 ;
      RECT 102.623 98.175 103.511 99.502 ;
      RECT 102.623 98.175 103.557 99.456 ;
      RECT 102.623 98.175 103.603 99.41 ;
      RECT 102.623 98.175 103.649 99.364 ;
      RECT 101.473 99.304 103.665 99.333 ;
      RECT 102.623 98.175 110 99.325 ;
      RECT 107.675 108.902 110 110 ;
      RECT 108.925 107.675 110 110 ;
      RECT 107.721 108.856 110 110 ;
      RECT 108.917 107.679 110 110 ;
      RECT 107.767 108.81 110 110 ;
      RECT 108.871 107.706 110 110 ;
      RECT 107.813 108.764 110 110 ;
      RECT 108.825 107.752 110 110 ;
      RECT 107.859 108.718 110 110 ;
      RECT 108.779 107.798 110 110 ;
      RECT 107.905 108.672 110 110 ;
      RECT 108.733 107.844 110 110 ;
      RECT 107.951 108.626 110 110 ;
      RECT 108.687 107.89 110 110 ;
      RECT 107.997 108.58 110 110 ;
      RECT 108.641 107.936 110 110 ;
      RECT 108.043 108.534 110 110 ;
      RECT 108.595 107.982 110 110 ;
      RECT 108.089 108.488 110 110 ;
      RECT 108.549 108.028 110 110 ;
      RECT 108.135 108.442 110 110 ;
      RECT 108.503 108.074 110 110 ;
      RECT 108.181 108.396 110 110 ;
      RECT 108.457 108.12 110 110 ;
      RECT 108.227 108.35 110 110 ;
      RECT 108.411 108.166 110 110 ;
      RECT 108.273 108.304 110 110 ;
      RECT 108.365 108.212 110 110 ;
      RECT 108.319 108.258 110 110 ;
    LAYER MET4 SPACING 0.1 ;
      RECT -20 -20 3.325 110 ;
      RECT -20 -20 3.371 55.817 ;
      RECT -20 -20 3.417 55.771 ;
      RECT -20 -20 3.463 55.725 ;
      RECT -20 -20 3.509 55.679 ;
      RECT -20 -20 3.555 55.633 ;
      RECT -20 -20 3.601 55.587 ;
      RECT -20 -20 3.647 55.541 ;
      RECT -20 -20 3.693 55.495 ;
      RECT -20 -20 3.739 55.449 ;
      RECT -20 -20 3.785 55.403 ;
      RECT -20 -20 3.831 55.357 ;
      RECT -20 -20 3.877 55.311 ;
      RECT -20 -20 3.923 55.265 ;
      RECT -20 -20 3.969 55.219 ;
      RECT -20 -20 4.015 55.173 ;
      RECT -20 -20 4.061 55.127 ;
      RECT -20 -20 4.107 55.081 ;
      RECT -20 -20 4.153 55.035 ;
      RECT -20 -20 4.199 54.989 ;
      RECT -20 -20 4.245 54.943 ;
      RECT -20 -20 4.291 54.897 ;
      RECT -20 -20 4.337 54.851 ;
      RECT -20 -20 4.383 54.805 ;
      RECT -20 -20 4.429 54.759 ;
      RECT -20 -20 4.475 54.713 ;
      RECT -20 -20 4.521 54.667 ;
      RECT -20 -20 4.567 54.621 ;
      RECT -20 -20 4.613 54.575 ;
      RECT -20 -20 4.659 54.529 ;
      RECT -20 -20 4.705 54.483 ;
      RECT -20 -20 4.751 54.437 ;
      RECT -20 -20 4.797 54.391 ;
      RECT -20 -20 4.843 54.345 ;
      RECT -20 -20 4.889 54.299 ;
      RECT -20 -20 4.935 54.253 ;
      RECT -20 -20 4.981 54.207 ;
      RECT -20 -20 5.027 54.161 ;
      RECT -20 -20 5.073 54.115 ;
      RECT -20 -20 5.119 54.069 ;
      RECT -20 -20 5.165 54.023 ;
      RECT -20 -20 5.211 53.977 ;
      RECT -20 -20 5.257 53.931 ;
      RECT -20 -20 5.303 53.885 ;
      RECT -20 -20 5.349 53.839 ;
      RECT -20 -20 5.395 53.793 ;
      RECT -20 -20 5.441 53.747 ;
      RECT -20 -20 5.487 53.701 ;
      RECT -20 -20 5.533 53.655 ;
      RECT -20 -20 5.579 53.609 ;
      RECT -20 -20 5.625 53.563 ;
      RECT -20 -20 5.671 53.517 ;
      RECT -20 -20 5.717 53.471 ;
      RECT -20 -20 5.763 53.425 ;
      RECT -20 -20 5.809 53.379 ;
      RECT -20 -20 5.855 53.333 ;
      RECT -20 -20 5.901 53.287 ;
      RECT -20 -20 5.947 53.241 ;
      RECT -20 -20 5.993 53.195 ;
      RECT -20 -20 6.039 53.149 ;
      RECT -20 -20 6.085 53.103 ;
      RECT -20 -20 6.131 53.057 ;
      RECT -20 -20 6.177 53.011 ;
      RECT -20 -20 6.223 52.965 ;
      RECT -20 -20 6.269 52.919 ;
      RECT -20 -20 6.315 52.873 ;
      RECT -20 -20 6.361 52.827 ;
      RECT -20 -20 6.407 52.781 ;
      RECT -20 -20 6.453 52.735 ;
      RECT -20 -20 6.499 52.689 ;
      RECT -20 -20 6.545 52.643 ;
      RECT -20 -20 6.591 52.597 ;
      RECT -20 -20 6.637 52.551 ;
      RECT -20 -20 6.683 52.505 ;
      RECT -20 -20 6.729 52.459 ;
      RECT -20 -20 6.775 52.413 ;
      RECT -20 -20 6.821 52.367 ;
      RECT -20 -20 6.867 52.321 ;
      RECT -20 -20 6.913 52.275 ;
      RECT -20 -20 6.959 52.229 ;
      RECT -20 -20 7.005 52.183 ;
      RECT -20 -20 7.051 52.137 ;
      RECT -20 -20 7.097 52.091 ;
      RECT -20 -20 7.143 52.045 ;
      RECT -20 -20 7.189 51.999 ;
      RECT -20 -20 7.235 51.953 ;
      RECT -20 -20 7.281 51.907 ;
      RECT -20 -20 7.327 51.861 ;
      RECT -20 -20 7.373 51.815 ;
      RECT -20 -20 7.419 51.769 ;
      RECT -20 -20 7.465 51.723 ;
      RECT -20 -20 7.511 51.677 ;
      RECT -20 -20 7.557 51.631 ;
      RECT -20 -20 7.603 51.585 ;
      RECT -20 -20 7.649 51.539 ;
      RECT -20 -20 7.695 51.493 ;
      RECT -20 -20 7.741 51.447 ;
      RECT -20 -20 7.787 51.401 ;
      RECT -20 -20 7.833 51.355 ;
      RECT -20 -20 7.879 51.309 ;
      RECT -20 -20 7.925 51.263 ;
      RECT -20 -20 7.971 51.217 ;
      RECT -20 -20 8.017 51.171 ;
      RECT -20 -20 8.063 51.125 ;
      RECT -20 -20 8.109 51.079 ;
      RECT -20 -20 8.155 51.033 ;
      RECT -20 -20 8.201 50.987 ;
      RECT -20 -20 8.247 50.941 ;
      RECT -20 -20 8.293 50.895 ;
      RECT -20 -20 8.339 50.849 ;
      RECT -20 -20 8.385 50.803 ;
      RECT -20 -20 8.431 50.757 ;
      RECT -20 -20 8.477 50.711 ;
      RECT -20 -20 8.523 50.665 ;
      RECT -20 -20 8.569 50.619 ;
      RECT -20 -20 8.615 50.573 ;
      RECT -20 -20 8.661 50.527 ;
      RECT -20 -20 8.707 50.481 ;
      RECT -20 -20 8.753 50.435 ;
      RECT -20 -20 8.799 50.389 ;
      RECT -20 -20 8.845 50.343 ;
      RECT -20 -20 8.891 50.297 ;
      RECT -20 -20 8.937 50.251 ;
      RECT -20 -20 8.983 50.205 ;
      RECT -20 -20 9.029 50.159 ;
      RECT -20 -20 9.075 50.113 ;
      RECT -20 -20 9.121 50.067 ;
      RECT -20 -20 9.167 50.021 ;
      RECT -20 -20 9.213 49.975 ;
      RECT -20 -20 9.259 49.929 ;
      RECT -20 -20 9.305 49.883 ;
      RECT -20 -20 9.351 49.837 ;
      RECT -20 -20 9.397 49.791 ;
      RECT -20 -20 9.443 49.745 ;
      RECT -20 -20 9.489 49.699 ;
      RECT -20 -20 9.535 49.653 ;
      RECT -20 -20 9.581 49.607 ;
      RECT -20 -20 9.627 49.561 ;
      RECT -20 -20 9.673 49.515 ;
      RECT -20 -20 9.719 49.469 ;
      RECT -20 -20 9.765 49.423 ;
      RECT -20 -20 9.811 49.377 ;
      RECT -20 -20 9.857 49.331 ;
      RECT -20 -20 9.903 49.285 ;
      RECT -20 -20 9.949 49.239 ;
      RECT -20 -20 9.995 49.193 ;
      RECT -20 -20 10.041 49.147 ;
      RECT -20 -20 10.087 49.101 ;
      RECT -20 -20 10.133 49.055 ;
      RECT -20 -20 10.179 49.009 ;
      RECT -20 -20 10.225 48.963 ;
      RECT -20 -20 10.271 48.917 ;
      RECT -20 -20 10.317 48.871 ;
      RECT -20 -20 10.363 48.825 ;
      RECT -20 -20 10.409 48.779 ;
      RECT -20 -20 10.455 48.733 ;
      RECT -20 -20 10.501 48.687 ;
      RECT -20 -20 10.547 48.641 ;
      RECT -20 -20 10.593 48.595 ;
      RECT -20 -20 10.639 48.549 ;
      RECT -20 -20 10.685 48.503 ;
      RECT -20 -20 10.731 48.457 ;
      RECT -20 -20 10.777 48.411 ;
      RECT -20 -20 10.823 48.365 ;
      RECT -20 -20 10.869 48.319 ;
      RECT -20 -20 10.915 48.273 ;
      RECT -20 -20 10.961 48.227 ;
      RECT -20 -20 11.007 48.181 ;
      RECT -20 -20 11.053 48.135 ;
      RECT -20 -20 11.099 48.089 ;
      RECT -20 -20 11.145 48.043 ;
      RECT -20 -20 11.191 47.997 ;
      RECT -20 -20 11.237 47.951 ;
      RECT -20 -20 11.283 47.905 ;
      RECT -20 -20 11.329 47.859 ;
      RECT -20 -20 11.375 47.813 ;
      RECT -20 -20 11.421 47.767 ;
      RECT -20 -20 11.467 47.721 ;
      RECT -20 -20 11.513 47.675 ;
      RECT -20 -20 11.559 47.629 ;
      RECT -20 -20 11.605 47.583 ;
      RECT -20 -20 11.651 47.537 ;
      RECT -20 -20 11.697 47.491 ;
      RECT -20 -20 11.743 47.445 ;
      RECT -20 -20 11.789 47.399 ;
      RECT -20 -20 11.835 47.353 ;
      RECT -20 -20 11.881 47.307 ;
      RECT -20 -20 11.927 47.261 ;
      RECT -20 -20 11.973 47.215 ;
      RECT -20 -20 12.019 47.169 ;
      RECT -20 -20 12.065 47.123 ;
      RECT -20 -20 12.111 47.077 ;
      RECT -20 -20 12.157 47.031 ;
      RECT -20 -20 12.203 46.985 ;
      RECT -20 -20 12.249 46.939 ;
      RECT -20 -20 12.295 46.893 ;
      RECT -20 -20 12.341 46.847 ;
      RECT -20 -20 12.387 46.801 ;
      RECT -20 -20 12.433 46.755 ;
      RECT -20 -20 12.479 46.709 ;
      RECT -20 -20 12.525 46.663 ;
      RECT -20 -20 12.571 46.617 ;
      RECT -20 -20 12.617 46.571 ;
      RECT -20 -20 12.663 46.525 ;
      RECT -20 -20 12.709 46.479 ;
      RECT -20 -20 12.755 46.433 ;
      RECT -20 -20 12.801 46.387 ;
      RECT -20 -20 12.847 46.341 ;
      RECT -20 -20 12.893 46.295 ;
      RECT -20 -20 12.939 46.249 ;
      RECT -20 -20 12.985 46.203 ;
      RECT -20 -20 13.031 46.157 ;
      RECT -20 -20 13.077 46.111 ;
      RECT -20 -20 13.123 46.065 ;
      RECT -20 -20 13.169 46.019 ;
      RECT -20 -20 13.215 45.973 ;
      RECT -20 -20 13.261 45.927 ;
      RECT -20 -20 13.307 45.881 ;
      RECT -20 -20 13.353 45.835 ;
      RECT -20 -20 13.399 45.789 ;
      RECT -20 -20 13.445 45.743 ;
      RECT -20 -20 13.491 45.697 ;
      RECT -20 -20 13.537 45.651 ;
      RECT -20 -20 13.583 45.605 ;
      RECT -20 -20 13.629 45.559 ;
      RECT -20 -20 13.675 45.513 ;
      RECT -20 -20 13.721 45.467 ;
      RECT -20 -20 13.767 45.421 ;
      RECT -20 -20 13.813 45.375 ;
      RECT -20 -20 13.859 45.329 ;
      RECT -20 -20 13.905 45.283 ;
      RECT -20 -20 13.951 45.237 ;
      RECT -20 -20 13.997 45.191 ;
      RECT -20 -20 14.043 45.145 ;
      RECT -20 -20 14.089 45.099 ;
      RECT -20 -20 14.135 45.053 ;
      RECT -20 -20 14.181 45.007 ;
      RECT -20 -20 14.227 44.961 ;
      RECT -20 -20 14.273 44.915 ;
      RECT -20 -20 14.319 44.869 ;
      RECT -20 -20 14.365 44.823 ;
      RECT -20 -20 14.411 44.777 ;
      RECT -20 -20 14.457 44.731 ;
      RECT -20 -20 14.503 44.685 ;
      RECT -20 -20 14.549 44.639 ;
      RECT -20 -20 14.595 44.593 ;
      RECT -20 -20 14.641 44.547 ;
      RECT -20 -20 14.687 44.501 ;
      RECT -20 -20 14.733 44.455 ;
      RECT -20 -20 14.779 44.409 ;
      RECT -20 -20 14.825 44.363 ;
      RECT -20 -20 14.871 44.317 ;
      RECT -20 -20 14.917 44.271 ;
      RECT -20 -20 14.963 44.225 ;
      RECT -20 -20 15.009 44.179 ;
      RECT -20 -20 15.055 44.133 ;
      RECT -20 -20 15.101 44.087 ;
      RECT -20 -20 15.147 44.041 ;
      RECT -20 -20 15.193 43.995 ;
      RECT -20 -20 15.239 43.949 ;
      RECT -20 -20 15.285 43.903 ;
      RECT -20 -20 15.325 43.86 ;
      RECT -20 -20 15.371 43.817 ;
      RECT -20 -20 15.417 43.771 ;
      RECT -20 -20 15.463 43.725 ;
      RECT -20 -20 15.509 43.679 ;
      RECT -20 -20 15.555 43.633 ;
      RECT -20 -20 15.601 43.587 ;
      RECT -20 -20 15.647 43.541 ;
      RECT -20 -20 15.693 43.495 ;
      RECT -20 -20 15.739 43.449 ;
      RECT -20 -20 15.785 43.403 ;
      RECT -20 -20 15.831 43.357 ;
      RECT -20 -20 15.877 43.311 ;
      RECT -20 -20 15.923 43.265 ;
      RECT -20 -20 15.969 43.219 ;
      RECT -20 -20 16.015 43.173 ;
      RECT -20 -20 16.061 43.127 ;
      RECT -20 -20 16.107 43.081 ;
      RECT -20 -20 16.153 43.035 ;
      RECT -20 -20 16.199 42.989 ;
      RECT -20 -20 16.245 42.943 ;
      RECT -20 -20 16.291 42.897 ;
      RECT -20 -20 16.337 42.851 ;
      RECT -20 -20 16.383 42.805 ;
      RECT -20 -20 16.429 42.759 ;
      RECT -20 -20 16.475 42.713 ;
      RECT -20 -20 16.521 42.667 ;
      RECT -20 -20 16.567 42.621 ;
      RECT -20 -20 16.613 42.575 ;
      RECT -20 -20 16.659 42.529 ;
      RECT -20 -20 16.705 42.483 ;
      RECT -20 -20 16.751 42.437 ;
      RECT -20 -20 16.797 42.391 ;
      RECT -20 -20 16.843 42.345 ;
      RECT -20 -20 16.889 42.299 ;
      RECT -20 -20 16.935 42.253 ;
      RECT -20 -20 16.981 42.207 ;
      RECT -20 -20 17.027 42.161 ;
      RECT -20 -20 17.073 42.115 ;
      RECT -20 -20 17.119 42.069 ;
      RECT -20 -20 17.165 42.023 ;
      RECT -20 -20 17.211 41.977 ;
      RECT -20 -20 17.257 41.931 ;
      RECT -20 -20 17.303 41.885 ;
      RECT -20 -20 17.349 41.839 ;
      RECT -20 -20 17.395 41.793 ;
      RECT -20 -20 17.441 41.747 ;
      RECT -20 -20 17.487 41.701 ;
      RECT -20 -20 17.533 41.655 ;
      RECT -20 -20 17.579 41.609 ;
      RECT -20 -20 17.625 41.563 ;
      RECT -20 -20 17.671 41.517 ;
      RECT -20 -20 17.717 41.471 ;
      RECT -20 -20 17.763 41.425 ;
      RECT -20 -20 17.809 41.379 ;
      RECT -20 -20 17.855 41.333 ;
      RECT -20 -20 17.901 41.287 ;
      RECT -20 -20 17.947 41.241 ;
      RECT -20 -20 17.993 41.195 ;
      RECT -20 -20 18.039 41.149 ;
      RECT -20 -20 18.085 41.103 ;
      RECT -20 -20 18.131 41.057 ;
      RECT -20 -20 18.177 41.011 ;
      RECT -20 -20 18.223 40.965 ;
      RECT -20 -20 18.269 40.919 ;
      RECT -20 -20 18.315 40.873 ;
      RECT -20 -20 18.361 40.827 ;
      RECT -20 -20 18.407 40.781 ;
      RECT -20 -20 18.453 40.735 ;
      RECT -20 -20 18.499 40.689 ;
      RECT -20 -20 18.545 40.643 ;
      RECT -20 -20 18.591 40.597 ;
      RECT -20 -20 18.637 40.551 ;
      RECT -20 -20 18.683 40.505 ;
      RECT -20 -20 18.729 40.459 ;
      RECT -20 -20 18.775 40.413 ;
      RECT -20 -20 18.821 40.367 ;
      RECT -20 -20 18.867 40.321 ;
      RECT -20 -20 18.913 40.275 ;
      RECT -20 -20 18.959 40.229 ;
      RECT -20 -20 19.005 40.183 ;
      RECT -20 -20 19.051 40.137 ;
      RECT -20 -20 19.097 40.091 ;
      RECT -20 -20 19.143 40.045 ;
      RECT -20 -20 19.189 39.999 ;
      RECT -20 -20 19.235 39.953 ;
      RECT -20 -20 19.281 39.907 ;
      RECT -20 -20 19.327 39.861 ;
      RECT -20 -20 19.373 39.815 ;
      RECT -20 -20 19.419 39.769 ;
      RECT -20 -20 19.465 39.723 ;
      RECT -20 -20 19.511 39.677 ;
      RECT -20 -20 19.557 39.631 ;
      RECT -20 -20 19.603 39.585 ;
      RECT -20 -20 19.649 39.539 ;
      RECT -20 -20 19.695 39.493 ;
      RECT -20 -20 19.741 39.447 ;
      RECT -20 -20 19.787 39.401 ;
      RECT -20 -20 19.833 39.355 ;
      RECT -20 -20 19.879 39.309 ;
      RECT -20 -20 19.925 39.263 ;
      RECT -20 -20 19.971 39.217 ;
      RECT -20 -20 20.017 39.171 ;
      RECT -20 -20 20.063 39.125 ;
      RECT -20 -20 20.109 39.079 ;
      RECT -20 -20 20.155 39.033 ;
      RECT -20 -20 20.201 38.987 ;
      RECT -20 -20 20.247 38.941 ;
      RECT -20 -20 20.293 38.895 ;
      RECT -20 -20 20.339 38.849 ;
      RECT -20 -20 20.385 38.803 ;
      RECT -20 -20 20.431 38.757 ;
      RECT -20 -20 20.477 38.711 ;
      RECT -20 -20 20.523 38.665 ;
      RECT -20 -20 20.569 38.619 ;
      RECT -20 -20 20.615 38.573 ;
      RECT -20 -20 20.661 38.527 ;
      RECT -20 -20 20.707 38.481 ;
      RECT -20 -20 20.753 38.435 ;
      RECT -20 -20 20.799 38.389 ;
      RECT -20 -20 20.845 38.343 ;
      RECT -20 -20 20.891 38.297 ;
      RECT -20 -20 20.937 38.251 ;
      RECT -20 -20 20.983 38.205 ;
      RECT -20 -20 21.029 38.159 ;
      RECT -20 -20 21.075 38.113 ;
      RECT -20 -20 21.121 38.067 ;
      RECT -20 -20 21.167 38.021 ;
      RECT -20 -20 21.213 37.975 ;
      RECT -20 -20 21.259 37.929 ;
      RECT -20 -20 21.305 37.883 ;
      RECT -20 -20 21.351 37.837 ;
      RECT -20 -20 21.397 37.791 ;
      RECT -20 -20 21.443 37.745 ;
      RECT -20 -20 21.489 37.699 ;
      RECT -20 -20 21.535 37.653 ;
      RECT -20 -20 21.581 37.607 ;
      RECT -20 -20 21.627 37.561 ;
      RECT -20 -20 21.673 37.515 ;
      RECT -20 -20 21.719 37.469 ;
      RECT -20 -20 21.765 37.423 ;
      RECT -20 -20 21.811 37.377 ;
      RECT -20 -20 21.857 37.331 ;
      RECT -20 -20 21.903 37.285 ;
      RECT -20 -20 21.949 37.239 ;
      RECT -20 -20 21.995 37.193 ;
      RECT -20 -20 22.041 37.147 ;
      RECT -20 -20 22.087 37.101 ;
      RECT -20 -20 22.133 37.055 ;
      RECT -20 -20 22.179 37.009 ;
      RECT -20 -20 22.225 36.963 ;
      RECT -20 -20 22.271 36.917 ;
      RECT -20 -20 22.317 36.871 ;
      RECT -20 -20 22.363 36.825 ;
      RECT -20 -20 22.409 36.779 ;
      RECT -20 -20 22.455 36.733 ;
      RECT -20 -20 22.501 36.687 ;
      RECT -20 -20 22.547 36.641 ;
      RECT -20 -20 22.593 36.595 ;
      RECT -20 -20 22.639 36.549 ;
      RECT -20 -20 22.685 36.503 ;
      RECT -20 -20 22.731 36.457 ;
      RECT -20 -20 22.777 36.411 ;
      RECT -20 -20 22.823 36.365 ;
      RECT -20 -20 22.869 36.319 ;
      RECT -20 -20 22.915 36.273 ;
      RECT -20 -20 22.961 36.227 ;
      RECT -20 -20 23.007 36.181 ;
      RECT -20 -20 23.053 36.135 ;
      RECT -20 -20 23.099 36.089 ;
      RECT -20 -20 23.145 36.043 ;
      RECT -20 -20 23.191 35.997 ;
      RECT -20 -20 23.237 35.951 ;
      RECT -20 -20 23.283 35.905 ;
      RECT -20 -20 23.329 35.859 ;
      RECT -20 -20 23.375 35.813 ;
      RECT -20 -20 23.421 35.767 ;
      RECT -20 -20 23.467 35.721 ;
      RECT -20 -20 23.513 35.675 ;
      RECT -20 -20 23.559 35.629 ;
      RECT -20 -20 23.605 35.583 ;
      RECT -20 -20 23.651 35.537 ;
      RECT -20 -20 23.697 35.491 ;
      RECT -20 -20 23.743 35.445 ;
      RECT -20 -20 23.789 35.399 ;
      RECT -20 -20 23.835 35.353 ;
      RECT -20 -20 23.881 35.307 ;
      RECT -20 -20 23.927 35.261 ;
      RECT -20 -20 23.973 35.215 ;
      RECT -20 -20 24.019 35.169 ;
      RECT -20 -20 24.065 35.123 ;
      RECT -20 -20 24.111 35.077 ;
      RECT -20 -20 24.157 35.031 ;
      RECT -20 -20 24.203 34.985 ;
      RECT -20 -20 24.249 34.939 ;
      RECT -20 -20 24.295 34.893 ;
      RECT -20 -20 24.341 34.847 ;
      RECT -20 -20 24.387 34.801 ;
      RECT -20 -20 24.433 34.755 ;
      RECT -20 -20 24.479 34.709 ;
      RECT -20 -20 24.525 34.663 ;
      RECT -20 -20 24.571 34.617 ;
      RECT -20 -20 24.617 34.571 ;
      RECT -20 -20 24.663 34.525 ;
      RECT -20 -20 24.709 34.479 ;
      RECT -20 -20 24.755 34.433 ;
      RECT -20 -20 24.801 34.387 ;
      RECT -20 -20 24.847 34.341 ;
      RECT -20 -20 24.893 34.295 ;
      RECT -20 -20 24.939 34.249 ;
      RECT -20 -20 24.985 34.203 ;
      RECT -20 -20 25.031 34.157 ;
      RECT -20 -20 25.077 34.111 ;
      RECT -20 -20 25.123 34.065 ;
      RECT -20 -20 25.169 34.019 ;
      RECT -20 -20 25.215 33.973 ;
      RECT -20 -20 25.261 33.927 ;
      RECT -20 -20 25.307 33.881 ;
      RECT -20 -20 25.353 33.835 ;
      RECT -20 -20 25.399 33.789 ;
      RECT -20 -20 25.445 33.743 ;
      RECT -20 -20 25.491 33.697 ;
      RECT -20 -20 25.537 33.651 ;
      RECT -20 -20 25.583 33.605 ;
      RECT -20 -20 25.629 33.559 ;
      RECT -20 -20 25.675 33.513 ;
      RECT -20 -20 25.721 33.467 ;
      RECT -20 -20 25.767 33.421 ;
      RECT -20 -20 25.813 33.375 ;
      RECT -20 -20 25.859 33.329 ;
      RECT -20 -20 25.905 33.283 ;
      RECT -20 -20 25.951 33.237 ;
      RECT -20 -20 25.997 33.191 ;
      RECT -20 -20 26.043 33.145 ;
      RECT -20 -20 26.089 33.099 ;
      RECT -20 -20 26.135 33.053 ;
      RECT -20 -20 26.181 33.007 ;
      RECT -20 -20 26.227 32.961 ;
      RECT -20 -20 26.273 32.915 ;
      RECT -20 -20 26.319 32.869 ;
      RECT -20 -20 26.365 32.823 ;
      RECT -20 -20 26.411 32.777 ;
      RECT -20 -20 26.457 32.731 ;
      RECT -20 -20 26.503 32.685 ;
      RECT -20 -20 26.549 32.639 ;
      RECT -20 -20 26.595 32.593 ;
      RECT -20 -20 26.641 32.547 ;
      RECT -20 -20 26.687 32.501 ;
      RECT -20 -20 26.733 32.455 ;
      RECT -20 -20 26.779 32.409 ;
      RECT -20 -20 26.825 32.363 ;
      RECT -20 -20 26.871 32.317 ;
      RECT -20 -20 26.917 32.271 ;
      RECT -20 -20 26.963 32.225 ;
      RECT -20 -20 27.009 32.179 ;
      RECT -20 -20 27.055 32.133 ;
      RECT -20 -20 27.101 32.087 ;
      RECT -20 -20 27.147 32.041 ;
      RECT -20 -20 27.193 31.995 ;
      RECT -20 -20 27.239 31.949 ;
      RECT -20 -20 27.285 31.903 ;
      RECT -20 -20 27.331 31.857 ;
      RECT -20 -20 27.377 31.811 ;
      RECT -20 -20 27.423 31.765 ;
      RECT -20 -20 27.469 31.719 ;
      RECT -20 -20 27.515 31.673 ;
      RECT -20 -20 27.561 31.627 ;
      RECT -20 -20 27.607 31.581 ;
      RECT -20 -20 27.653 31.535 ;
      RECT -20 -20 27.699 31.489 ;
      RECT -20 -20 27.745 31.443 ;
      RECT -20 -20 27.791 31.397 ;
      RECT -20 -20 27.837 31.351 ;
      RECT -20 -20 27.883 31.305 ;
      RECT -20 -20 27.929 31.259 ;
      RECT -20 -20 27.975 31.213 ;
      RECT -20 -20 28.021 31.167 ;
      RECT -20 -20 28.067 31.121 ;
      RECT -20 -20 28.113 31.075 ;
      RECT -20 -20 28.159 31.029 ;
      RECT -20 -20 28.205 30.983 ;
      RECT -20 -20 28.251 30.937 ;
      RECT -20 -20 28.297 30.891 ;
      RECT -20 -20 28.343 30.845 ;
      RECT -20 -20 28.389 30.799 ;
      RECT -20 -20 28.435 30.753 ;
      RECT -20 -20 28.481 30.707 ;
      RECT -20 -20 28.527 30.661 ;
      RECT -20 -20 28.573 30.615 ;
      RECT -20 -20 28.619 30.569 ;
      RECT -20 -20 28.665 30.523 ;
      RECT -20 -20 28.711 30.477 ;
      RECT -20 -20 28.757 30.431 ;
      RECT -20 -20 28.803 30.385 ;
      RECT -20 -20 28.849 30.339 ;
      RECT -20 -20 28.895 30.293 ;
      RECT -20 -20 28.941 30.247 ;
      RECT -20 -20 28.987 30.201 ;
      RECT -20 -20 29.033 30.155 ;
      RECT -20 -20 29.079 30.109 ;
      RECT -20 -20 29.125 30.063 ;
      RECT -20 -20 29.171 30.017 ;
      RECT -20 -20 29.217 29.971 ;
      RECT -20 -20 29.263 29.925 ;
      RECT -20 -20 29.309 29.879 ;
      RECT -20 -20 29.355 29.833 ;
      RECT -20 -20 29.401 29.787 ;
      RECT -20 -20 29.447 29.741 ;
      RECT -20 -20 29.493 29.695 ;
      RECT -20 -20 29.539 29.649 ;
      RECT -20 -20 29.585 29.603 ;
      RECT -20 -20 29.631 29.557 ;
      RECT -20 -20 29.677 29.511 ;
      RECT -20 -20 29.723 29.465 ;
      RECT -20 -20 29.769 29.419 ;
      RECT -20 -20 29.815 29.373 ;
      RECT -20 -20 29.861 29.327 ;
      RECT -20 -20 29.907 29.281 ;
      RECT -20 -20 29.953 29.235 ;
      RECT -20 -20 29.999 29.189 ;
      RECT -20 -20 30.045 29.143 ;
      RECT -20 -20 30.091 29.097 ;
      RECT -20 -20 30.137 29.051 ;
      RECT -20 -20 30.183 29.005 ;
      RECT -20 -20 30.229 28.959 ;
      RECT -20 -20 30.275 28.913 ;
      RECT -20 -20 30.321 28.867 ;
      RECT -20 -20 30.367 28.821 ;
      RECT -20 -20 30.413 28.775 ;
      RECT -20 -20 30.459 28.729 ;
      RECT -20 -20 30.505 28.683 ;
      RECT -20 -20 30.551 28.637 ;
      RECT -20 -20 30.597 28.591 ;
      RECT -20 -20 30.643 28.545 ;
      RECT -20 -20 30.689 28.499 ;
      RECT -20 -20 30.735 28.453 ;
      RECT -20 -20 30.781 28.407 ;
      RECT -20 -20 30.827 28.361 ;
      RECT -20 -20 30.873 28.315 ;
      RECT -20 -20 30.919 28.269 ;
      RECT -20 -20 30.965 28.223 ;
      RECT -20 -20 31.011 28.177 ;
      RECT -20 -20 31.057 28.131 ;
      RECT -20 -20 31.103 28.085 ;
      RECT -20 -20 31.149 28.039 ;
      RECT -20 -20 31.195 27.993 ;
      RECT -20 -20 31.241 27.947 ;
      RECT -20 -20 31.287 27.901 ;
      RECT -20 -20 31.333 27.855 ;
      RECT -20 -20 31.379 27.809 ;
      RECT -20 -20 31.425 27.763 ;
      RECT -20 -20 31.471 27.717 ;
      RECT -20 -20 31.517 27.671 ;
      RECT -20 -20 31.563 27.625 ;
      RECT -20 -20 31.609 27.579 ;
      RECT -20 -20 31.655 27.533 ;
      RECT -20 -20 31.701 27.487 ;
      RECT -20 -20 31.747 27.441 ;
      RECT -20 -20 31.793 27.395 ;
      RECT -20 -20 31.839 27.349 ;
      RECT -20 -20 31.885 27.303 ;
      RECT -20 -20 31.931 27.257 ;
      RECT -20 -20 31.977 27.211 ;
      RECT -20 -20 32.023 27.165 ;
      RECT -20 -20 32.069 27.119 ;
      RECT -20 -20 32.115 27.073 ;
      RECT -20 -20 32.161 27.027 ;
      RECT -20 -20 32.207 26.981 ;
      RECT -20 -20 32.253 26.935 ;
      RECT -20 -20 32.299 26.889 ;
      RECT -20 -20 32.345 26.843 ;
      RECT -20 -20 32.391 26.797 ;
      RECT -20 -20 32.437 26.751 ;
      RECT -20 -20 32.483 26.705 ;
      RECT -20 -20 32.529 26.659 ;
      RECT -20 -20 32.575 26.613 ;
      RECT -20 -20 32.621 26.567 ;
      RECT -20 -20 32.667 26.521 ;
      RECT -20 -20 32.713 26.475 ;
      RECT -20 -20 32.759 26.429 ;
      RECT -20 -20 32.805 26.383 ;
      RECT -20 -20 32.851 26.337 ;
      RECT -20 -20 32.897 26.291 ;
      RECT -20 -20 32.943 26.245 ;
      RECT -20 -20 32.989 26.199 ;
      RECT -20 -20 33.035 26.153 ;
      RECT -20 -20 33.081 26.107 ;
      RECT -20 -20 33.127 26.061 ;
      RECT -20 -20 33.173 26.015 ;
      RECT -20 -20 33.219 25.969 ;
      RECT -20 -20 33.265 25.923 ;
      RECT -20 -20 33.311 25.877 ;
      RECT -20 -20 33.357 25.831 ;
      RECT -20 -20 33.403 25.785 ;
      RECT -20 -20 33.449 25.739 ;
      RECT -20 -20 33.495 25.693 ;
      RECT -20 -20 33.541 25.647 ;
      RECT -20 -20 33.587 25.601 ;
      RECT -20 -20 33.633 25.555 ;
      RECT -20 -20 33.679 25.509 ;
      RECT -20 -20 33.725 25.463 ;
      RECT -20 -20 33.771 25.417 ;
      RECT -20 -20 33.817 25.371 ;
      RECT -20 -20 33.863 25.325 ;
      RECT -20 -20 33.909 25.279 ;
      RECT -20 -20 33.955 25.233 ;
      RECT -20 -20 34.001 25.187 ;
      RECT -20 -20 34.047 25.141 ;
      RECT -20 -20 34.093 25.095 ;
      RECT -20 -20 34.139 25.049 ;
      RECT -20 -20 34.185 25.003 ;
      RECT -20 -20 34.231 24.957 ;
      RECT -20 -20 34.277 24.911 ;
      RECT -20 -20 34.323 24.865 ;
      RECT -20 -20 34.369 24.819 ;
      RECT -20 -20 34.415 24.773 ;
      RECT -20 -20 34.461 24.727 ;
      RECT -20 -20 34.507 24.681 ;
      RECT -20 -20 34.553 24.635 ;
      RECT -20 -20 34.599 24.589 ;
      RECT -20 -20 34.645 24.543 ;
      RECT -20 -20 34.691 24.497 ;
      RECT -20 -20 34.737 24.451 ;
      RECT -20 -20 34.783 24.405 ;
      RECT -20 -20 34.829 24.359 ;
      RECT -20 -20 34.875 24.313 ;
      RECT -20 -20 34.921 24.267 ;
      RECT -20 -20 34.967 24.221 ;
      RECT -20 -20 35.013 24.175 ;
      RECT -20 -20 35.059 24.129 ;
      RECT -20 -20 35.105 24.083 ;
      RECT -20 -20 35.151 24.037 ;
      RECT -20 -20 35.197 23.991 ;
      RECT -20 -20 35.243 23.945 ;
      RECT -20 -20 35.289 23.899 ;
      RECT -20 -20 35.335 23.853 ;
      RECT -20 -20 35.381 23.807 ;
      RECT -20 -20 35.427 23.761 ;
      RECT -20 -20 35.473 23.715 ;
      RECT -20 -20 35.519 23.669 ;
      RECT -20 -20 35.565 23.623 ;
      RECT -20 -20 35.611 23.577 ;
      RECT -20 -20 35.657 23.531 ;
      RECT -20 -20 35.703 23.485 ;
      RECT -20 -20 35.749 23.439 ;
      RECT -20 -20 35.795 23.393 ;
      RECT -20 -20 35.841 23.347 ;
      RECT -20 -20 35.887 23.301 ;
      RECT -20 -20 35.933 23.255 ;
      RECT -20 -20 35.979 23.209 ;
      RECT -20 -20 36.025 23.163 ;
      RECT -20 -20 36.071 23.117 ;
      RECT -20 -20 36.117 23.071 ;
      RECT -20 -20 36.163 23.025 ;
      RECT -20 -20 36.209 22.979 ;
      RECT -20 -20 36.255 22.933 ;
      RECT -20 -20 36.301 22.887 ;
      RECT -20 -20 36.347 22.841 ;
      RECT -20 -20 36.393 22.795 ;
      RECT -20 -20 36.439 22.749 ;
      RECT -20 -20 36.485 22.703 ;
      RECT -20 -20 36.531 22.657 ;
      RECT -20 -20 36.577 22.611 ;
      RECT -20 -20 36.623 22.565 ;
      RECT -20 -20 36.669 22.519 ;
      RECT -20 -20 36.715 22.473 ;
      RECT -20 -20 36.761 22.427 ;
      RECT -20 -20 36.807 22.381 ;
      RECT -20 -20 36.853 22.335 ;
      RECT -20 -20 36.899 22.289 ;
      RECT -20 -20 36.945 22.243 ;
      RECT -20 -20 36.991 22.197 ;
      RECT -20 -20 37.037 22.151 ;
      RECT -20 -20 37.083 22.105 ;
      RECT -20 -20 37.129 22.059 ;
      RECT -20 -20 37.175 22.013 ;
      RECT -20 -20 37.221 21.967 ;
      RECT -20 -20 37.267 21.921 ;
      RECT -20 -20 37.313 21.875 ;
      RECT -20 -20 37.359 21.829 ;
      RECT -20 -20 37.405 21.783 ;
      RECT -20 -20 37.451 21.737 ;
      RECT -20 -20 37.497 21.691 ;
      RECT -20 -20 37.543 21.645 ;
      RECT -20 -20 37.589 21.599 ;
      RECT -20 -20 37.635 21.553 ;
      RECT -20 -20 37.681 21.507 ;
      RECT -20 -20 37.727 21.461 ;
      RECT -20 -20 37.773 21.415 ;
      RECT -20 -20 37.819 21.369 ;
      RECT -20 -20 37.865 21.323 ;
      RECT -20 -20 37.911 21.277 ;
      RECT -20 -20 37.957 21.231 ;
      RECT -20 -20 38.003 21.185 ;
      RECT -20 -20 38.049 21.139 ;
      RECT -20 -20 38.095 21.093 ;
      RECT -20 -20 38.141 21.047 ;
      RECT -20 -20 38.187 21.001 ;
      RECT -20 -20 38.233 20.955 ;
      RECT -20 -20 38.279 20.909 ;
      RECT -20 -20 38.325 20.863 ;
      RECT -20 -20 38.371 20.817 ;
      RECT -20 -20 38.417 20.771 ;
      RECT -20 -20 38.463 20.725 ;
      RECT -20 -20 38.509 20.679 ;
      RECT -20 -20 38.555 20.633 ;
      RECT -20 -20 38.601 20.587 ;
      RECT -20 -20 38.647 20.541 ;
      RECT -20 -20 38.693 20.495 ;
      RECT -20 -20 38.739 20.449 ;
      RECT -20 -20 38.785 20.403 ;
      RECT -20 -20 38.831 20.357 ;
      RECT -20 -20 38.877 20.311 ;
      RECT -20 -20 38.923 20.265 ;
      RECT -20 -20 38.969 20.219 ;
      RECT -20 -20 39.015 20.173 ;
      RECT -20 -20 39.061 20.127 ;
      RECT -20 -20 39.107 20.081 ;
      RECT -20 -20 39.153 20.035 ;
      RECT -20 -20 39.199 19.989 ;
      RECT -20 -20 39.245 19.943 ;
      RECT -20 -20 39.291 19.897 ;
      RECT -20 -20 39.337 19.851 ;
      RECT -20 -20 39.383 19.805 ;
      RECT -20 -20 39.429 19.759 ;
      RECT -20 -20 39.475 19.713 ;
      RECT -20 -20 39.521 19.667 ;
      RECT -20 -20 39.567 19.621 ;
      RECT -20 -20 39.613 19.575 ;
      RECT -20 -20 39.659 19.529 ;
      RECT -20 -20 39.705 19.483 ;
      RECT -20 -20 39.751 19.437 ;
      RECT -20 -20 39.797 19.391 ;
      RECT -20 -20 39.843 19.345 ;
      RECT -20 -20 39.889 19.299 ;
      RECT -20 -20 39.935 19.253 ;
      RECT -20 -20 39.981 19.207 ;
      RECT -20 -20 40.027 19.161 ;
      RECT -20 -20 40.073 19.115 ;
      RECT -20 -20 40.119 19.069 ;
      RECT -20 -20 40.165 19.023 ;
      RECT -20 -20 40.211 18.977 ;
      RECT -20 -20 40.257 18.931 ;
      RECT -20 -20 40.303 18.885 ;
      RECT -20 -20 40.349 18.839 ;
      RECT -20 -20 40.395 18.793 ;
      RECT -20 -20 40.441 18.747 ;
      RECT -20 -20 40.487 18.701 ;
      RECT -20 -20 40.533 18.655 ;
      RECT -20 -20 40.579 18.609 ;
      RECT -20 -20 40.625 18.563 ;
      RECT -20 -20 40.671 18.517 ;
      RECT -20 -20 40.717 18.471 ;
      RECT -20 -20 40.763 18.425 ;
      RECT -20 -20 40.809 18.379 ;
      RECT -20 -20 40.855 18.333 ;
      RECT -20 -20 40.901 18.287 ;
      RECT -20 -20 40.947 18.241 ;
      RECT -20 -20 40.993 18.195 ;
      RECT -20 -20 41.039 18.149 ;
      RECT -20 -20 41.085 18.103 ;
      RECT -20 -20 41.131 18.057 ;
      RECT -20 -20 41.177 18.011 ;
      RECT -20 -20 41.223 17.965 ;
      RECT -20 -20 41.269 17.919 ;
      RECT -20 -20 41.315 17.873 ;
      RECT -20 -20 41.361 17.827 ;
      RECT -20 -20 41.407 17.781 ;
      RECT -20 -20 41.453 17.735 ;
      RECT -20 -20 41.499 17.689 ;
      RECT -20 -20 41.545 17.643 ;
      RECT -20 -20 41.591 17.597 ;
      RECT -20 -20 41.637 17.551 ;
      RECT -20 -20 41.683 17.505 ;
      RECT -20 -20 41.729 17.459 ;
      RECT -20 -20 41.775 17.413 ;
      RECT -20 -20 41.821 17.367 ;
      RECT -20 -20 41.867 17.321 ;
      RECT -20 -20 41.913 17.275 ;
      RECT -20 -20 41.959 17.229 ;
      RECT -20 -20 42.005 17.183 ;
      RECT -20 -20 42.051 17.137 ;
      RECT -20 -20 42.097 17.091 ;
      RECT -20 -20 42.143 17.045 ;
      RECT -20 -20 42.189 16.999 ;
      RECT -20 -20 42.235 16.953 ;
      RECT -20 -20 42.281 16.907 ;
      RECT -20 -20 42.327 16.861 ;
      RECT -20 -20 42.373 16.815 ;
      RECT -20 -20 42.419 16.769 ;
      RECT -20 -20 42.465 16.723 ;
      RECT -20 -20 42.511 16.677 ;
      RECT -20 -20 42.557 16.631 ;
      RECT -20 -20 42.603 16.585 ;
      RECT -20 -20 42.649 16.539 ;
      RECT -20 -20 42.695 16.493 ;
      RECT -20 -20 42.741 16.447 ;
      RECT -20 -20 42.787 16.401 ;
      RECT -20 -20 42.833 16.355 ;
      RECT -20 -20 42.879 16.309 ;
      RECT -20 -20 42.925 16.263 ;
      RECT -20 -20 42.971 16.217 ;
      RECT -20 -20 43.017 16.171 ;
      RECT -20 -20 43.063 16.125 ;
      RECT -20 -20 43.109 16.079 ;
      RECT -20 -20 43.155 16.033 ;
      RECT -20 -20 43.201 15.987 ;
      RECT -20 -20 43.247 15.941 ;
      RECT -20 -20 43.293 15.895 ;
      RECT -20 -20 43.339 15.849 ;
      RECT -20 -20 43.385 15.803 ;
      RECT -20 -20 43.431 15.757 ;
      RECT -20 -20 43.477 15.711 ;
      RECT -20 -20 43.523 15.665 ;
      RECT -20 -20 43.569 15.619 ;
      RECT -20 -20 43.615 15.573 ;
      RECT -20 -20 43.661 15.527 ;
      RECT -20 -20 43.707 15.481 ;
      RECT -20 -20 43.753 15.435 ;
      RECT -20 -20 43.799 15.389 ;
      RECT -20 -20 43.845 15.343 ;
      RECT -20 -20 43.891 15.297 ;
      RECT -20 -20 43.937 15.251 ;
      RECT -20 -20 43.983 15.205 ;
      RECT -20 -20 44.029 15.159 ;
      RECT -20 -20 44.075 15.113 ;
      RECT -20 -20 44.121 15.067 ;
      RECT -20 -20 44.167 15.021 ;
      RECT -20 -20 44.213 14.975 ;
      RECT -20 -20 44.259 14.929 ;
      RECT -20 -20 44.305 14.883 ;
      RECT -20 -20 44.351 14.837 ;
      RECT -20 -20 44.397 14.791 ;
      RECT -20 -20 44.443 14.745 ;
      RECT -20 -20 44.489 14.699 ;
      RECT -20 -20 44.535 14.653 ;
      RECT -20 -20 44.581 14.607 ;
      RECT -20 -20 44.627 14.561 ;
      RECT -20 -20 44.673 14.515 ;
      RECT -20 -20 44.719 14.469 ;
      RECT -20 -20 44.765 14.423 ;
      RECT -20 -20 44.811 14.377 ;
      RECT -20 -20 44.857 14.331 ;
      RECT -20 -20 44.903 14.285 ;
      RECT -20 -20 44.949 14.239 ;
      RECT -20 -20 44.995 14.193 ;
      RECT -20 -20 45.041 14.147 ;
      RECT -20 -20 45.087 14.101 ;
      RECT -20 -20 45.133 14.055 ;
      RECT -20 -20 45.179 14.009 ;
      RECT -20 -20 45.225 13.963 ;
      RECT -20 -20 45.271 13.917 ;
      RECT -20 -20 45.317 13.871 ;
      RECT -20 -20 45.363 13.825 ;
      RECT -20 -20 45.409 13.779 ;
      RECT -20 -20 45.455 13.733 ;
      RECT -20 -20 45.501 13.687 ;
      RECT -20 -20 45.547 13.641 ;
      RECT -20 -20 45.593 13.595 ;
      RECT -20 -20 45.639 13.549 ;
      RECT -20 -20 45.685 13.503 ;
      RECT -20 -20 45.731 13.457 ;
      RECT -20 -20 45.777 13.411 ;
      RECT -20 -20 45.823 13.365 ;
      RECT -20 -20 45.869 13.319 ;
      RECT -20 -20 45.915 13.273 ;
      RECT -20 -20 45.961 13.227 ;
      RECT -20 -20 46.007 13.181 ;
      RECT -20 -20 46.053 13.135 ;
      RECT -20 -20 46.099 13.089 ;
      RECT -20 -20 46.145 13.043 ;
      RECT -20 -20 46.191 12.997 ;
      RECT -20 -20 46.237 12.951 ;
      RECT -20 -20 46.283 12.905 ;
      RECT -20 -20 46.329 12.859 ;
      RECT -20 -20 46.375 12.813 ;
      RECT -20 -20 46.421 12.767 ;
      RECT -20 -20 46.467 12.721 ;
      RECT -20 -20 46.513 12.675 ;
      RECT -20 -20 46.559 12.629 ;
      RECT -20 -20 46.605 12.583 ;
      RECT -20 -20 46.651 12.537 ;
      RECT -20 -20 46.697 12.491 ;
      RECT -20 -20 46.743 12.445 ;
      RECT -20 -20 46.789 12.399 ;
      RECT -20 -20 46.835 12.353 ;
      RECT -20 -20 46.881 12.307 ;
      RECT -20 -20 46.927 12.261 ;
      RECT -20 -20 46.973 12.215 ;
      RECT -20 -20 47.019 12.169 ;
      RECT -20 -20 47.065 12.123 ;
      RECT -20 -20 47.111 12.077 ;
      RECT -20 -20 47.157 12.031 ;
      RECT -20 -20 47.203 11.985 ;
      RECT -20 -20 47.249 11.939 ;
      RECT -20 -20 47.295 11.893 ;
      RECT -20 -20 47.341 11.847 ;
      RECT -20 -20 47.387 11.801 ;
      RECT -20 -20 47.433 11.755 ;
      RECT -20 -20 47.479 11.709 ;
      RECT -20 -20 47.525 11.663 ;
      RECT -20 -20 47.571 11.617 ;
      RECT -20 -20 47.617 11.571 ;
      RECT -20 -20 47.663 11.525 ;
      RECT -20 -20 47.709 11.479 ;
      RECT -20 -20 47.755 11.433 ;
      RECT -20 -20 47.801 11.387 ;
      RECT -20 -20 47.847 11.341 ;
      RECT -20 -20 47.893 11.295 ;
      RECT -20 -20 47.939 11.249 ;
      RECT -20 -20 47.985 11.203 ;
      RECT -20 -20 48.031 11.157 ;
      RECT -20 -20 48.077 11.111 ;
      RECT -20 -20 48.123 11.065 ;
      RECT -20 -20 48.169 11.019 ;
      RECT -20 -20 48.215 10.973 ;
      RECT -20 -20 48.261 10.927 ;
      RECT -20 -20 48.307 10.881 ;
      RECT -20 -20 48.353 10.835 ;
      RECT -20 -20 48.399 10.789 ;
      RECT -20 -20 48.445 10.743 ;
      RECT -20 -20 48.491 10.697 ;
      RECT -20 -20 48.537 10.651 ;
      RECT -20 -20 48.583 10.605 ;
      RECT -20 -20 48.629 10.559 ;
      RECT -20 -20 48.675 10.513 ;
      RECT -20 -20 48.721 10.467 ;
      RECT -20 -20 48.767 10.421 ;
      RECT -20 -20 48.813 10.375 ;
      RECT -20 -20 48.859 10.329 ;
      RECT -20 -20 48.905 10.283 ;
      RECT -20 -20 48.951 10.237 ;
      RECT -20 -20 48.997 10.191 ;
      RECT -20 -20 49.043 10.145 ;
      RECT -20 -20 49.089 10.099 ;
      RECT -20 -20 49.135 10.053 ;
      RECT -20 -20 49.181 10.007 ;
      RECT -20 -20 49.227 9.961 ;
      RECT -20 -20 49.273 9.915 ;
      RECT -20 -20 49.319 9.869 ;
      RECT -20 -20 49.365 9.823 ;
      RECT -20 -20 49.411 9.777 ;
      RECT -20 -20 49.457 9.731 ;
      RECT -20 -20 49.503 9.685 ;
      RECT -20 -20 49.549 9.639 ;
      RECT -20 -20 49.595 9.593 ;
      RECT -20 -20 49.641 9.547 ;
      RECT -20 -20 49.687 9.501 ;
      RECT -20 -20 49.733 9.455 ;
      RECT -20 -20 49.779 9.409 ;
      RECT -20 -20 49.825 9.363 ;
      RECT -20 -20 49.871 9.317 ;
      RECT -20 -20 49.917 9.271 ;
      RECT -20 -20 49.963 9.225 ;
      RECT -20 -20 50.009 9.179 ;
      RECT -20 -20 50.055 9.133 ;
      RECT -20 -20 50.101 9.087 ;
      RECT -20 -20 50.147 9.041 ;
      RECT -20 -20 50.193 8.995 ;
      RECT -20 -20 50.239 8.949 ;
      RECT -20 -20 50.285 8.903 ;
      RECT -20 -20 50.331 8.857 ;
      RECT -20 -20 50.377 8.811 ;
      RECT -20 -20 50.423 8.765 ;
      RECT -20 -20 50.469 8.719 ;
      RECT -20 -20 50.515 8.673 ;
      RECT -20 -20 50.561 8.627 ;
      RECT -20 -20 50.607 8.581 ;
      RECT -20 -20 50.653 8.535 ;
      RECT -20 -20 50.699 8.489 ;
      RECT -20 -20 50.745 8.443 ;
      RECT -20 -20 50.791 8.397 ;
      RECT -20 -20 50.837 8.351 ;
      RECT -20 -20 50.883 8.305 ;
      RECT -20 -20 50.929 8.259 ;
      RECT -20 -20 50.975 8.213 ;
      RECT -20 -20 51.021 8.167 ;
      RECT -20 -20 51.067 8.121 ;
      RECT -20 -20 51.113 8.075 ;
      RECT -20 -20 51.159 8.029 ;
      RECT -20 -20 51.205 7.983 ;
      RECT -20 -20 51.251 7.937 ;
      RECT -20 -20 51.297 7.891 ;
      RECT -20 -20 51.343 7.845 ;
      RECT -20 -20 51.389 7.799 ;
      RECT -20 -20 51.435 7.753 ;
      RECT -20 -20 51.481 7.707 ;
      RECT -20 -20 51.527 7.661 ;
      RECT -20 -20 51.573 7.615 ;
      RECT -20 -20 51.619 7.569 ;
      RECT -20 -20 51.665 7.523 ;
      RECT -20 -20 51.711 7.477 ;
      RECT -20 -20 51.757 7.431 ;
      RECT -20 -20 51.803 7.385 ;
      RECT -20 -20 51.849 7.339 ;
      RECT -20 -20 51.895 7.293 ;
      RECT -20 -20 51.941 7.247 ;
      RECT -20 -20 51.987 7.201 ;
      RECT -20 -20 52.033 7.155 ;
      RECT -20 -20 52.079 7.109 ;
      RECT -20 -20 52.125 7.063 ;
      RECT -20 -20 52.171 7.017 ;
      RECT -20 -20 52.217 6.971 ;
      RECT -20 -20 52.263 6.925 ;
      RECT -20 -20 52.309 6.879 ;
      RECT -20 -20 52.355 6.833 ;
      RECT -20 -20 52.401 6.787 ;
      RECT -20 -20 52.447 6.741 ;
      RECT -20 -20 52.493 6.695 ;
      RECT -20 -20 52.539 6.649 ;
      RECT -20 -20 52.585 6.603 ;
      RECT -20 -20 52.631 6.557 ;
      RECT -20 -20 52.677 6.511 ;
      RECT -20 -20 52.723 6.465 ;
      RECT -20 -20 52.769 6.419 ;
      RECT -20 -20 52.815 6.373 ;
      RECT -20 -20 52.861 6.327 ;
      RECT -20 -20 52.907 6.281 ;
      RECT -20 -20 52.953 6.235 ;
      RECT -20 -20 52.999 6.189 ;
      RECT -20 -20 53.045 6.143 ;
      RECT -20 -20 53.091 6.097 ;
      RECT -20 -20 53.137 6.051 ;
      RECT -20 -20 53.183 6.005 ;
      RECT -20 -20 53.229 5.959 ;
      RECT -20 -20 53.275 5.913 ;
      RECT -20 -20 53.321 5.867 ;
      RECT -20 -20 53.367 5.821 ;
      RECT -20 -20 53.413 5.775 ;
      RECT -20 -20 53.459 5.729 ;
      RECT -20 -20 53.505 5.683 ;
      RECT -20 -20 53.551 5.637 ;
      RECT -20 -20 53.597 5.591 ;
      RECT -20 -20 53.643 5.545 ;
      RECT -20 -20 53.689 5.499 ;
      RECT -20 -20 53.735 5.453 ;
      RECT -20 -20 53.781 5.407 ;
      RECT -20 -20 53.827 5.361 ;
      RECT -20 -20 53.873 5.315 ;
      RECT -20 -20 53.919 5.269 ;
      RECT -20 -20 53.965 5.223 ;
      RECT -20 -20 54.011 5.177 ;
      RECT -20 -20 54.057 5.131 ;
      RECT -20 -20 54.103 5.085 ;
      RECT -20 -20 54.149 5.039 ;
      RECT -20 -20 54.195 4.993 ;
      RECT -20 -20 54.241 4.947 ;
      RECT -20 -20 54.287 4.901 ;
      RECT -20 -20 54.333 4.855 ;
      RECT -20 -20 54.379 4.809 ;
      RECT -20 -20 54.425 4.763 ;
      RECT -20 -20 54.471 4.717 ;
      RECT -20 -20 54.517 4.671 ;
      RECT -20 -20 54.563 4.625 ;
      RECT -20 -20 54.609 4.579 ;
      RECT -20 -20 54.655 4.533 ;
      RECT -20 -20 54.701 4.487 ;
      RECT -20 -20 54.747 4.441 ;
      RECT -20 -20 54.793 4.395 ;
      RECT -20 -20 54.839 4.349 ;
      RECT -20 -20 54.885 4.303 ;
      RECT -20 -20 54.931 4.257 ;
      RECT -20 -20 54.977 4.211 ;
      RECT -20 -20 55.023 4.165 ;
      RECT -20 -20 55.069 4.119 ;
      RECT -20 -20 55.115 4.073 ;
      RECT -20 -20 55.161 4.027 ;
      RECT -20 -20 55.207 3.981 ;
      RECT -20 -20 55.253 3.935 ;
      RECT -20 -20 55.299 3.889 ;
      RECT -20 -20 55.345 3.843 ;
      RECT -20 -20 55.391 3.797 ;
      RECT -20 -20 55.437 3.751 ;
      RECT -20 -20 55.483 3.705 ;
      RECT -20 -20 55.529 3.659 ;
      RECT -20 -20 55.575 3.613 ;
      RECT -20 -20 55.621 3.567 ;
      RECT -20 -20 55.667 3.521 ;
      RECT -20 -20 55.713 3.475 ;
      RECT -20 -20 55.759 3.429 ;
      RECT -20 -20 55.805 3.383 ;
      RECT -20 -20 55.84 3.342 ;
      RECT -20 -20 110 3.325 ;
      RECT 15.675 61.137 16.825 110 ;
      RECT 15.675 61.137 16.871 62.567 ;
      RECT 15.675 61.137 16.917 62.521 ;
      RECT 15.675 61.137 16.963 62.475 ;
      RECT 15.675 61.137 17.009 62.429 ;
      RECT 15.675 61.137 17.055 62.383 ;
      RECT 15.675 61.137 17.101 62.337 ;
      RECT 15.675 61.137 17.147 62.291 ;
      RECT 15.675 61.137 17.193 62.245 ;
      RECT 15.675 61.137 17.239 62.199 ;
      RECT 15.675 61.137 17.285 62.153 ;
      RECT 15.675 61.137 17.331 62.107 ;
      RECT 15.675 61.137 17.377 62.061 ;
      RECT 15.675 61.137 17.423 62.015 ;
      RECT 15.675 61.137 17.469 61.969 ;
      RECT 15.675 61.137 17.515 61.923 ;
      RECT 15.675 61.137 17.561 61.877 ;
      RECT 15.675 61.137 17.607 61.831 ;
      RECT 15.675 61.137 17.653 61.785 ;
      RECT 15.675 61.137 17.699 61.739 ;
      RECT 15.675 61.137 17.745 61.693 ;
      RECT 15.675 61.137 17.791 61.647 ;
      RECT 15.675 61.137 17.837 61.601 ;
      RECT 15.675 61.137 17.883 61.555 ;
      RECT 15.675 61.137 17.929 61.509 ;
      RECT 15.675 61.137 17.975 61.463 ;
      RECT 15.675 61.137 18.021 61.417 ;
      RECT 15.675 61.137 18.067 61.371 ;
      RECT 15.675 61.137 18.113 61.325 ;
      RECT 15.675 61.137 18.159 61.279 ;
      RECT 15.675 61.137 18.205 61.233 ;
      RECT 15.675 61.137 18.251 61.187 ;
      RECT 15.721 61.091 18.297 61.141 ;
      RECT 15.767 61.045 18.343 61.095 ;
      RECT 15.813 60.999 18.389 61.049 ;
      RECT 15.859 60.953 18.435 61.003 ;
      RECT 15.905 60.907 18.481 60.957 ;
      RECT 15.951 60.861 18.527 60.911 ;
      RECT 15.997 60.815 18.573 60.865 ;
      RECT 16.043 60.769 18.619 60.819 ;
      RECT 16.089 60.723 18.665 60.773 ;
      RECT 16.135 60.677 18.711 60.727 ;
      RECT 16.181 60.631 18.757 60.681 ;
      RECT 16.227 60.585 18.803 60.635 ;
      RECT 16.273 60.539 18.849 60.589 ;
      RECT 16.319 60.493 18.895 60.543 ;
      RECT 16.365 60.447 18.941 60.497 ;
      RECT 16.411 60.401 18.987 60.451 ;
      RECT 16.457 60.355 19.033 60.405 ;
      RECT 16.503 60.309 19.079 60.359 ;
      RECT 16.549 60.263 19.125 60.313 ;
      RECT 16.595 60.217 19.171 60.267 ;
      RECT 16.641 60.171 19.217 60.221 ;
      RECT 16.687 60.125 19.263 60.175 ;
      RECT 16.733 60.079 19.309 60.129 ;
      RECT 16.779 60.033 19.355 60.083 ;
      RECT 16.825 59.987 19.401 60.037 ;
      RECT 16.871 59.941 19.447 59.991 ;
      RECT 16.917 59.895 19.493 59.945 ;
      RECT 16.963 59.849 19.539 59.899 ;
      RECT 17.009 59.803 19.585 59.853 ;
      RECT 17.055 59.757 19.631 59.807 ;
      RECT 17.101 59.711 19.677 59.761 ;
      RECT 17.147 59.665 19.723 59.715 ;
      RECT 17.193 59.619 19.769 59.669 ;
      RECT 17.239 59.573 19.815 59.623 ;
      RECT 17.285 59.527 19.861 59.577 ;
      RECT 17.331 59.481 19.907 59.531 ;
      RECT 17.377 59.435 19.953 59.485 ;
      RECT 17.423 59.389 19.999 59.439 ;
      RECT 17.469 59.343 20.045 59.393 ;
      RECT 17.515 59.297 20.091 59.347 ;
      RECT 17.561 59.251 20.137 59.301 ;
      RECT 17.607 59.205 20.183 59.255 ;
      RECT 17.653 59.159 20.229 59.209 ;
      RECT 17.699 59.113 20.275 59.163 ;
      RECT 17.745 59.067 20.321 59.117 ;
      RECT 17.791 59.021 20.367 59.071 ;
      RECT 17.837 58.975 20.413 59.025 ;
      RECT 17.883 58.929 20.459 58.979 ;
      RECT 17.929 58.883 20.505 58.933 ;
      RECT 17.975 58.837 20.551 58.887 ;
      RECT 18.021 58.791 20.597 58.841 ;
      RECT 18.067 58.745 20.643 58.795 ;
      RECT 18.113 58.699 20.689 58.749 ;
      RECT 18.159 58.653 20.735 58.703 ;
      RECT 18.205 58.607 20.781 58.657 ;
      RECT 18.251 58.561 20.827 58.611 ;
      RECT 18.297 58.515 20.873 58.565 ;
      RECT 18.343 58.469 20.919 58.519 ;
      RECT 18.389 58.423 20.965 58.473 ;
      RECT 18.435 58.377 21.011 58.427 ;
      RECT 18.481 58.331 21.057 58.381 ;
      RECT 18.527 58.285 21.103 58.335 ;
      RECT 18.573 58.239 21.149 58.289 ;
      RECT 18.619 58.193 21.195 58.243 ;
      RECT 18.665 58.147 21.241 58.197 ;
      RECT 18.711 58.101 21.287 58.151 ;
      RECT 18.757 58.055 21.333 58.105 ;
      RECT 18.803 58.009 21.379 58.059 ;
      RECT 18.849 57.963 21.425 58.013 ;
      RECT 18.895 57.917 21.471 57.967 ;
      RECT 18.941 57.871 21.517 57.921 ;
      RECT 18.987 57.825 21.563 57.875 ;
      RECT 19.033 57.779 21.609 57.829 ;
      RECT 19.079 57.733 21.655 57.783 ;
      RECT 19.125 57.687 21.701 57.737 ;
      RECT 19.171 57.641 21.747 57.691 ;
      RECT 19.217 57.595 21.793 57.645 ;
      RECT 19.263 57.549 21.839 57.599 ;
      RECT 19.309 57.503 21.885 57.553 ;
      RECT 19.355 57.457 21.931 57.507 ;
      RECT 19.401 57.411 21.977 57.461 ;
      RECT 19.447 57.365 22.023 57.415 ;
      RECT 19.493 57.319 22.069 57.369 ;
      RECT 19.539 57.273 22.115 57.323 ;
      RECT 19.585 57.227 22.161 57.277 ;
      RECT 19.631 57.181 22.207 57.231 ;
      RECT 19.677 57.135 22.253 57.185 ;
      RECT 19.723 57.089 22.299 57.139 ;
      RECT 19.769 57.043 22.345 57.093 ;
      RECT 19.815 56.997 22.391 57.047 ;
      RECT 19.861 56.951 22.437 57.001 ;
      RECT 19.907 56.905 22.483 56.955 ;
      RECT 19.953 56.859 22.529 56.909 ;
      RECT 19.999 56.813 22.575 56.863 ;
      RECT 20.045 56.767 22.621 56.817 ;
      RECT 20.091 56.721 22.667 56.771 ;
      RECT 20.137 56.675 22.713 56.725 ;
      RECT 20.183 56.629 22.759 56.679 ;
      RECT 20.229 56.583 22.805 56.633 ;
      RECT 20.275 56.537 22.851 56.587 ;
      RECT 20.321 56.491 22.897 56.541 ;
      RECT 20.367 56.445 22.943 56.495 ;
      RECT 20.413 56.399 22.989 56.449 ;
      RECT 20.459 56.353 23.035 56.403 ;
      RECT 20.505 56.307 23.081 56.357 ;
      RECT 20.551 56.261 23.127 56.311 ;
      RECT 20.597 56.215 23.173 56.265 ;
      RECT 20.643 56.169 23.219 56.219 ;
      RECT 20.689 56.123 23.265 56.173 ;
      RECT 20.735 56.077 23.311 56.127 ;
      RECT 20.781 56.031 23.357 56.081 ;
      RECT 20.827 55.985 23.403 56.035 ;
      RECT 20.873 55.939 23.449 55.989 ;
      RECT 20.919 55.893 23.495 55.943 ;
      RECT 20.965 55.847 23.541 55.897 ;
      RECT 21.011 55.801 23.587 55.851 ;
      RECT 21.057 55.755 23.633 55.805 ;
      RECT 21.103 55.709 23.679 55.759 ;
      RECT 21.149 55.663 23.725 55.713 ;
      RECT 21.195 55.617 23.771 55.667 ;
      RECT 21.241 55.571 23.817 55.621 ;
      RECT 21.287 55.525 23.863 55.575 ;
      RECT 21.333 55.479 23.909 55.529 ;
      RECT 21.379 55.433 23.955 55.483 ;
      RECT 21.425 55.387 24.001 55.437 ;
      RECT 21.471 55.341 24.047 55.391 ;
      RECT 21.517 55.295 24.093 55.345 ;
      RECT 21.563 55.249 24.139 55.299 ;
      RECT 21.609 55.203 24.185 55.253 ;
      RECT 21.655 55.157 24.231 55.207 ;
      RECT 21.701 55.111 24.277 55.161 ;
      RECT 21.747 55.065 24.323 55.115 ;
      RECT 21.793 55.019 24.369 55.069 ;
      RECT 21.839 54.973 24.415 55.023 ;
      RECT 21.885 54.927 24.461 54.977 ;
      RECT 21.931 54.881 24.507 54.931 ;
      RECT 21.977 54.835 24.553 54.885 ;
      RECT 22.023 54.789 24.599 54.839 ;
      RECT 22.069 54.743 24.645 54.793 ;
      RECT 22.115 54.697 24.691 54.747 ;
      RECT 22.161 54.651 24.737 54.701 ;
      RECT 22.207 54.605 24.783 54.655 ;
      RECT 22.253 54.559 24.829 54.609 ;
      RECT 22.299 54.513 24.875 54.563 ;
      RECT 22.345 54.467 24.921 54.517 ;
      RECT 22.391 54.421 24.967 54.471 ;
      RECT 22.437 54.375 25.013 54.425 ;
      RECT 22.483 54.329 25.059 54.379 ;
      RECT 22.529 54.283 25.105 54.333 ;
      RECT 22.575 54.237 25.151 54.287 ;
      RECT 22.621 54.191 25.197 54.241 ;
      RECT 22.667 54.145 25.243 54.195 ;
      RECT 22.713 54.099 25.289 54.149 ;
      RECT 22.759 54.053 25.335 54.103 ;
      RECT 22.805 54.007 25.381 54.057 ;
      RECT 22.851 53.961 25.427 54.011 ;
      RECT 22.897 53.915 25.473 53.965 ;
      RECT 22.943 53.869 25.519 53.919 ;
      RECT 22.989 53.823 25.565 53.873 ;
      RECT 23.035 53.777 25.611 53.827 ;
      RECT 23.081 53.731 25.657 53.781 ;
      RECT 23.127 53.685 25.703 53.735 ;
      RECT 23.173 53.639 25.749 53.689 ;
      RECT 23.219 53.593 25.795 53.643 ;
      RECT 23.265 53.547 25.841 53.597 ;
      RECT 23.311 53.501 25.887 53.551 ;
      RECT 23.357 53.455 25.933 53.505 ;
      RECT 23.403 53.409 25.979 53.459 ;
      RECT 23.449 53.363 26.025 53.413 ;
      RECT 23.495 53.317 26.071 53.367 ;
      RECT 23.541 53.271 26.117 53.321 ;
      RECT 23.587 53.225 26.163 53.275 ;
      RECT 23.633 53.179 26.209 53.229 ;
      RECT 23.679 53.133 26.255 53.183 ;
      RECT 23.725 53.087 26.301 53.137 ;
      RECT 23.771 53.041 26.347 53.091 ;
      RECT 23.817 52.995 26.393 53.045 ;
      RECT 23.863 52.949 26.439 52.999 ;
      RECT 23.909 52.903 26.485 52.953 ;
      RECT 23.955 52.857 26.531 52.907 ;
      RECT 24.001 52.811 26.577 52.861 ;
      RECT 24.047 52.765 26.623 52.815 ;
      RECT 24.093 52.719 26.669 52.769 ;
      RECT 24.139 52.673 26.715 52.723 ;
      RECT 24.185 52.627 26.761 52.677 ;
      RECT 24.231 52.581 26.807 52.631 ;
      RECT 24.277 52.535 26.853 52.585 ;
      RECT 24.323 52.489 26.899 52.539 ;
      RECT 24.369 52.443 26.945 52.493 ;
      RECT 24.415 52.397 26.991 52.447 ;
      RECT 24.461 52.351 27.037 52.401 ;
      RECT 24.507 52.305 27.083 52.355 ;
      RECT 24.553 52.259 27.129 52.309 ;
      RECT 24.599 52.213 27.175 52.263 ;
      RECT 24.645 52.167 27.221 52.217 ;
      RECT 24.691 52.121 27.267 52.171 ;
      RECT 24.737 52.075 27.313 52.125 ;
      RECT 24.783 52.029 27.359 52.079 ;
      RECT 24.829 51.983 27.405 52.033 ;
      RECT 24.875 51.937 27.451 51.987 ;
      RECT 24.921 51.891 27.497 51.941 ;
      RECT 24.967 51.845 27.543 51.895 ;
      RECT 25.013 51.799 27.589 51.849 ;
      RECT 25.059 51.753 27.635 51.803 ;
      RECT 25.105 51.707 27.681 51.757 ;
      RECT 25.151 51.661 27.727 51.711 ;
      RECT 25.197 51.615 27.773 51.665 ;
      RECT 25.243 51.569 27.819 51.619 ;
      RECT 25.289 51.523 27.865 51.573 ;
      RECT 25.335 51.477 27.911 51.527 ;
      RECT 25.381 51.431 27.957 51.481 ;
      RECT 25.427 51.385 28.003 51.435 ;
      RECT 25.473 51.339 28.049 51.389 ;
      RECT 25.519 51.293 28.095 51.343 ;
      RECT 25.565 51.247 28.141 51.297 ;
      RECT 25.611 51.201 28.187 51.251 ;
      RECT 25.657 51.155 28.233 51.205 ;
      RECT 25.703 51.109 28.279 51.159 ;
      RECT 25.749 51.063 28.325 51.113 ;
      RECT 25.795 51.017 28.371 51.067 ;
      RECT 25.841 50.971 28.417 51.021 ;
      RECT 25.887 50.925 28.463 50.975 ;
      RECT 25.933 50.879 28.509 50.929 ;
      RECT 25.979 50.833 28.555 50.883 ;
      RECT 26.025 50.787 28.601 50.837 ;
      RECT 26.071 50.741 28.647 50.791 ;
      RECT 26.117 50.695 28.693 50.745 ;
      RECT 26.163 50.649 28.739 50.699 ;
      RECT 26.209 50.603 28.785 50.653 ;
      RECT 26.255 50.557 28.825 50.61 ;
      RECT 26.301 50.511 28.871 50.567 ;
      RECT 26.347 50.465 28.917 50.521 ;
      RECT 26.393 50.419 28.963 50.475 ;
      RECT 26.439 50.373 29.009 50.429 ;
      RECT 26.485 50.327 29.055 50.383 ;
      RECT 26.531 50.281 29.101 50.337 ;
      RECT 26.577 50.235 29.147 50.291 ;
      RECT 26.623 50.189 29.193 50.245 ;
      RECT 26.669 50.143 29.239 50.199 ;
      RECT 26.715 50.097 29.285 50.153 ;
      RECT 26.761 50.051 29.331 50.107 ;
      RECT 26.807 50.005 29.377 50.061 ;
      RECT 26.853 49.959 29.423 50.015 ;
      RECT 26.899 49.913 29.469 49.969 ;
      RECT 26.945 49.867 29.515 49.923 ;
      RECT 26.991 49.821 29.561 49.877 ;
      RECT 27.037 49.775 29.607 49.831 ;
      RECT 27.083 49.729 29.653 49.785 ;
      RECT 27.129 49.683 29.699 49.739 ;
      RECT 27.175 49.637 29.745 49.693 ;
      RECT 27.221 49.591 29.791 49.647 ;
      RECT 27.267 49.545 29.837 49.601 ;
      RECT 27.313 49.499 29.883 49.555 ;
      RECT 27.359 49.453 29.929 49.509 ;
      RECT 27.405 49.407 29.975 49.463 ;
      RECT 27.451 49.361 30.021 49.417 ;
      RECT 27.497 49.315 30.067 49.371 ;
      RECT 27.543 49.269 30.113 49.325 ;
      RECT 27.589 49.223 30.159 49.279 ;
      RECT 27.635 49.177 30.205 49.233 ;
      RECT 27.681 49.131 30.251 49.187 ;
      RECT 27.727 49.085 30.297 49.141 ;
      RECT 27.773 49.039 30.343 49.095 ;
      RECT 27.819 48.993 30.389 49.049 ;
      RECT 27.865 48.947 30.435 49.003 ;
      RECT 27.911 48.901 30.481 48.957 ;
      RECT 27.957 48.855 30.527 48.911 ;
      RECT 28.003 48.809 30.573 48.865 ;
      RECT 28.049 48.763 30.619 48.819 ;
      RECT 28.095 48.717 30.665 48.773 ;
      RECT 28.141 48.671 30.711 48.727 ;
      RECT 28.187 48.625 30.757 48.681 ;
      RECT 28.233 48.579 30.803 48.635 ;
      RECT 28.279 48.533 30.849 48.589 ;
      RECT 28.325 48.487 30.895 48.543 ;
      RECT 28.371 48.441 30.941 48.497 ;
      RECT 28.417 48.395 30.987 48.451 ;
      RECT 28.463 48.349 31.033 48.405 ;
      RECT 28.509 48.303 31.079 48.359 ;
      RECT 28.555 48.257 31.125 48.313 ;
      RECT 28.601 48.211 31.171 48.267 ;
      RECT 28.647 48.165 31.217 48.221 ;
      RECT 28.693 48.119 31.263 48.175 ;
      RECT 28.739 48.073 31.309 48.129 ;
      RECT 28.785 48.027 31.355 48.083 ;
      RECT 28.831 47.981 31.401 48.037 ;
      RECT 28.877 47.935 31.447 47.991 ;
      RECT 28.923 47.889 31.493 47.945 ;
      RECT 28.969 47.843 31.539 47.899 ;
      RECT 29.015 47.797 31.585 47.853 ;
      RECT 29.061 47.751 31.631 47.807 ;
      RECT 29.107 47.705 31.677 47.761 ;
      RECT 29.153 47.659 31.723 47.715 ;
      RECT 29.199 47.613 31.769 47.669 ;
      RECT 29.245 47.567 31.815 47.623 ;
      RECT 29.291 47.521 31.861 47.577 ;
      RECT 29.337 47.475 31.907 47.531 ;
      RECT 29.383 47.429 31.953 47.485 ;
      RECT 29.429 47.383 31.999 47.439 ;
      RECT 29.475 47.337 32.045 47.393 ;
      RECT 29.521 47.291 32.091 47.347 ;
      RECT 29.567 47.245 32.137 47.301 ;
      RECT 29.613 47.199 32.183 47.255 ;
      RECT 29.659 47.153 32.229 47.209 ;
      RECT 29.705 47.107 32.275 47.163 ;
      RECT 29.751 47.061 32.321 47.117 ;
      RECT 29.797 47.015 32.367 47.071 ;
      RECT 29.843 46.969 32.413 47.025 ;
      RECT 29.889 46.923 32.459 46.979 ;
      RECT 29.935 46.877 32.505 46.933 ;
      RECT 29.981 46.831 32.551 46.887 ;
      RECT 30.027 46.785 32.597 46.841 ;
      RECT 30.073 46.739 32.643 46.795 ;
      RECT 30.119 46.693 32.689 46.749 ;
      RECT 30.165 46.647 32.735 46.703 ;
      RECT 30.211 46.601 32.781 46.657 ;
      RECT 30.257 46.555 32.827 46.611 ;
      RECT 30.303 46.509 32.873 46.565 ;
      RECT 30.349 46.463 32.919 46.519 ;
      RECT 30.395 46.417 32.965 46.473 ;
      RECT 30.441 46.371 33.011 46.427 ;
      RECT 30.487 46.325 33.057 46.381 ;
      RECT 30.533 46.279 33.103 46.335 ;
      RECT 30.579 46.233 33.149 46.289 ;
      RECT 30.625 46.187 33.195 46.243 ;
      RECT 30.671 46.141 33.241 46.197 ;
      RECT 30.717 46.095 33.287 46.151 ;
      RECT 30.763 46.049 33.333 46.105 ;
      RECT 30.809 46.003 33.379 46.059 ;
      RECT 30.855 45.957 33.425 46.013 ;
      RECT 30.901 45.911 33.471 45.967 ;
      RECT 30.947 45.865 33.517 45.921 ;
      RECT 30.993 45.819 33.563 45.875 ;
      RECT 31.039 45.773 33.609 45.829 ;
      RECT 31.085 45.727 33.655 45.783 ;
      RECT 31.131 45.681 33.701 45.737 ;
      RECT 31.177 45.635 33.747 45.691 ;
      RECT 31.223 45.589 33.793 45.645 ;
      RECT 31.269 45.543 33.839 45.599 ;
      RECT 31.315 45.497 33.885 45.553 ;
      RECT 31.361 45.451 33.931 45.507 ;
      RECT 31.407 45.405 33.977 45.461 ;
      RECT 31.453 45.359 34.023 45.415 ;
      RECT 31.499 45.313 34.069 45.369 ;
      RECT 31.545 45.267 34.115 45.323 ;
      RECT 31.591 45.221 34.161 45.277 ;
      RECT 31.637 45.175 34.207 45.231 ;
      RECT 31.683 45.129 34.253 45.185 ;
      RECT 31.729 45.083 34.299 45.139 ;
      RECT 31.775 45.037 34.345 45.093 ;
      RECT 31.821 44.991 34.391 45.047 ;
      RECT 31.867 44.945 34.437 45.001 ;
      RECT 31.913 44.899 34.483 44.955 ;
      RECT 31.959 44.853 34.529 44.909 ;
      RECT 32.005 44.807 34.575 44.863 ;
      RECT 32.051 44.761 34.621 44.817 ;
      RECT 32.097 44.715 34.667 44.771 ;
      RECT 32.143 44.669 34.713 44.725 ;
      RECT 32.189 44.623 34.759 44.679 ;
      RECT 32.235 44.577 34.805 44.633 ;
      RECT 32.281 44.531 34.851 44.587 ;
      RECT 32.327 44.485 34.897 44.541 ;
      RECT 32.373 44.439 34.943 44.495 ;
      RECT 32.419 44.393 34.989 44.449 ;
      RECT 32.465 44.347 35.035 44.403 ;
      RECT 32.511 44.301 35.081 44.357 ;
      RECT 32.557 44.255 35.127 44.311 ;
      RECT 32.603 44.209 35.173 44.265 ;
      RECT 32.649 44.163 35.219 44.219 ;
      RECT 32.695 44.117 35.265 44.173 ;
      RECT 32.741 44.071 35.311 44.127 ;
      RECT 32.787 44.025 35.357 44.081 ;
      RECT 32.833 43.979 35.403 44.035 ;
      RECT 32.879 43.933 35.449 43.989 ;
      RECT 32.925 43.887 35.495 43.943 ;
      RECT 32.971 43.841 35.541 43.897 ;
      RECT 33.017 43.795 35.587 43.851 ;
      RECT 33.063 43.749 35.633 43.805 ;
      RECT 33.109 43.703 35.679 43.759 ;
      RECT 33.155 43.657 35.725 43.713 ;
      RECT 33.201 43.611 35.771 43.667 ;
      RECT 33.247 43.565 35.817 43.621 ;
      RECT 33.293 43.519 35.863 43.575 ;
      RECT 33.339 43.473 35.909 43.529 ;
      RECT 33.385 43.427 35.955 43.483 ;
      RECT 33.431 43.381 36.001 43.437 ;
      RECT 33.477 43.335 36.047 43.391 ;
      RECT 33.523 43.289 36.093 43.345 ;
      RECT 33.569 43.243 36.139 43.299 ;
      RECT 33.615 43.197 36.185 43.253 ;
      RECT 33.661 43.151 36.231 43.207 ;
      RECT 33.707 43.105 36.277 43.161 ;
      RECT 33.753 43.059 36.323 43.115 ;
      RECT 33.799 43.013 36.369 43.069 ;
      RECT 33.845 42.967 36.415 43.023 ;
      RECT 33.891 42.921 36.461 42.977 ;
      RECT 33.937 42.875 36.507 42.931 ;
      RECT 33.983 42.829 36.553 42.885 ;
      RECT 34.029 42.783 36.599 42.839 ;
      RECT 34.075 42.737 36.645 42.793 ;
      RECT 34.121 42.691 36.691 42.747 ;
      RECT 34.167 42.645 36.737 42.701 ;
      RECT 34.213 42.599 36.783 42.655 ;
      RECT 34.259 42.553 36.829 42.609 ;
      RECT 34.305 42.507 36.875 42.563 ;
      RECT 34.351 42.461 36.921 42.517 ;
      RECT 34.397 42.415 36.967 42.471 ;
      RECT 34.443 42.369 37.013 42.425 ;
      RECT 34.489 42.323 37.059 42.379 ;
      RECT 34.535 42.277 37.105 42.333 ;
      RECT 34.581 42.231 37.151 42.287 ;
      RECT 34.627 42.185 37.197 42.241 ;
      RECT 34.673 42.139 37.243 42.195 ;
      RECT 34.719 42.093 37.289 42.149 ;
      RECT 34.765 42.047 37.335 42.103 ;
      RECT 34.811 42.001 37.381 42.057 ;
      RECT 34.857 41.955 37.427 42.011 ;
      RECT 34.903 41.909 37.473 41.965 ;
      RECT 34.949 41.863 37.519 41.919 ;
      RECT 34.995 41.817 37.565 41.873 ;
      RECT 35.041 41.771 37.611 41.827 ;
      RECT 35.087 41.725 37.657 41.781 ;
      RECT 35.133 41.679 37.703 41.735 ;
      RECT 35.179 41.633 37.749 41.689 ;
      RECT 35.225 41.587 37.795 41.643 ;
      RECT 35.271 41.541 37.841 41.597 ;
      RECT 35.317 41.495 37.887 41.551 ;
      RECT 35.363 41.449 37.933 41.505 ;
      RECT 35.409 41.403 37.979 41.459 ;
      RECT 35.455 41.357 38.025 41.413 ;
      RECT 35.501 41.311 38.071 41.367 ;
      RECT 35.547 41.265 38.117 41.321 ;
      RECT 35.593 41.219 38.163 41.275 ;
      RECT 35.639 41.173 38.209 41.229 ;
      RECT 35.685 41.127 38.255 41.183 ;
      RECT 35.731 41.081 38.301 41.137 ;
      RECT 35.777 41.035 38.347 41.091 ;
      RECT 35.823 40.989 38.393 41.045 ;
      RECT 35.869 40.943 38.439 40.999 ;
      RECT 35.915 40.897 38.485 40.953 ;
      RECT 35.961 40.851 38.531 40.907 ;
      RECT 36.007 40.805 38.577 40.861 ;
      RECT 36.053 40.759 38.623 40.815 ;
      RECT 36.099 40.713 38.669 40.769 ;
      RECT 36.145 40.667 38.715 40.723 ;
      RECT 36.191 40.621 38.761 40.677 ;
      RECT 36.237 40.575 38.807 40.631 ;
      RECT 36.283 40.529 38.853 40.585 ;
      RECT 36.329 40.483 38.899 40.539 ;
      RECT 36.375 40.437 38.945 40.493 ;
      RECT 36.421 40.391 38.991 40.447 ;
      RECT 36.467 40.345 39.037 40.401 ;
      RECT 36.513 40.299 39.083 40.355 ;
      RECT 36.559 40.253 39.129 40.309 ;
      RECT 36.605 40.207 39.175 40.263 ;
      RECT 36.651 40.161 39.221 40.217 ;
      RECT 36.697 40.115 39.267 40.171 ;
      RECT 36.743 40.069 39.313 40.125 ;
      RECT 36.789 40.023 39.359 40.079 ;
      RECT 36.835 39.977 39.405 40.033 ;
      RECT 36.881 39.931 39.451 39.987 ;
      RECT 36.927 39.885 39.497 39.941 ;
      RECT 36.973 39.839 39.543 39.895 ;
      RECT 37.019 39.793 39.589 39.849 ;
      RECT 37.065 39.747 39.635 39.803 ;
      RECT 37.111 39.701 39.681 39.757 ;
      RECT 37.157 39.655 39.727 39.711 ;
      RECT 37.203 39.609 39.773 39.665 ;
      RECT 37.249 39.563 39.819 39.619 ;
      RECT 37.295 39.517 39.865 39.573 ;
      RECT 37.341 39.471 39.911 39.527 ;
      RECT 37.387 39.425 39.957 39.481 ;
      RECT 37.433 39.379 40.003 39.435 ;
      RECT 37.479 39.333 40.049 39.389 ;
      RECT 37.525 39.287 40.095 39.343 ;
      RECT 37.571 39.241 40.141 39.297 ;
      RECT 37.617 39.195 40.187 39.251 ;
      RECT 37.663 39.149 40.233 39.205 ;
      RECT 37.709 39.103 40.279 39.159 ;
      RECT 37.755 39.057 40.325 39.113 ;
      RECT 37.801 39.011 40.371 39.067 ;
      RECT 37.847 38.965 40.417 39.021 ;
      RECT 37.893 38.919 40.463 38.975 ;
      RECT 37.939 38.873 40.509 38.929 ;
      RECT 37.985 38.827 40.555 38.883 ;
      RECT 38.031 38.781 40.601 38.837 ;
      RECT 38.077 38.735 40.647 38.791 ;
      RECT 38.123 38.689 40.693 38.745 ;
      RECT 38.169 38.643 40.739 38.699 ;
      RECT 38.215 38.597 40.785 38.653 ;
      RECT 38.261 38.551 40.831 38.607 ;
      RECT 38.307 38.505 40.877 38.561 ;
      RECT 38.353 38.459 40.923 38.515 ;
      RECT 38.399 38.413 40.969 38.469 ;
      RECT 38.445 38.367 41.015 38.423 ;
      RECT 38.491 38.321 41.061 38.377 ;
      RECT 38.537 38.275 41.107 38.331 ;
      RECT 38.583 38.229 41.153 38.285 ;
      RECT 38.629 38.183 41.199 38.239 ;
      RECT 38.675 38.137 41.245 38.193 ;
      RECT 38.721 38.091 41.291 38.147 ;
      RECT 38.767 38.045 41.337 38.101 ;
      RECT 38.813 37.999 41.383 38.055 ;
      RECT 38.859 37.953 41.429 38.009 ;
      RECT 38.905 37.907 41.475 37.963 ;
      RECT 38.951 37.861 41.521 37.917 ;
      RECT 38.997 37.815 41.567 37.871 ;
      RECT 39.043 37.769 41.613 37.825 ;
      RECT 39.089 37.723 41.659 37.779 ;
      RECT 39.135 37.677 41.705 37.733 ;
      RECT 39.181 37.631 41.751 37.687 ;
      RECT 39.227 37.585 41.797 37.641 ;
      RECT 39.273 37.539 41.843 37.595 ;
      RECT 39.319 37.493 41.889 37.549 ;
      RECT 39.365 37.447 41.935 37.503 ;
      RECT 39.411 37.401 41.981 37.457 ;
      RECT 39.457 37.355 42.027 37.411 ;
      RECT 39.503 37.309 42.073 37.365 ;
      RECT 39.549 37.263 42.119 37.319 ;
      RECT 39.595 37.217 42.165 37.273 ;
      RECT 39.641 37.171 42.211 37.227 ;
      RECT 39.687 37.125 42.257 37.181 ;
      RECT 39.733 37.079 42.303 37.135 ;
      RECT 39.779 37.033 42.349 37.089 ;
      RECT 39.825 36.987 42.395 37.043 ;
      RECT 39.871 36.941 42.441 36.997 ;
      RECT 39.917 36.895 42.487 36.951 ;
      RECT 39.963 36.849 42.533 36.905 ;
      RECT 40.009 36.803 42.579 36.859 ;
      RECT 40.055 36.757 42.625 36.813 ;
      RECT 40.101 36.711 42.671 36.767 ;
      RECT 40.147 36.665 42.717 36.721 ;
      RECT 40.193 36.619 42.763 36.675 ;
      RECT 40.239 36.573 42.809 36.629 ;
      RECT 40.285 36.527 42.855 36.583 ;
      RECT 40.331 36.481 42.901 36.537 ;
      RECT 40.377 36.435 42.947 36.491 ;
      RECT 40.423 36.389 42.993 36.445 ;
      RECT 40.469 36.343 43.039 36.399 ;
      RECT 40.515 36.297 43.085 36.353 ;
      RECT 40.561 36.251 43.131 36.307 ;
      RECT 40.607 36.205 43.177 36.261 ;
      RECT 40.653 36.159 43.223 36.215 ;
      RECT 40.699 36.113 43.269 36.169 ;
      RECT 40.745 36.067 43.315 36.123 ;
      RECT 40.791 36.021 43.361 36.077 ;
      RECT 40.837 35.975 43.407 36.031 ;
      RECT 40.883 35.929 43.453 35.985 ;
      RECT 40.929 35.883 43.499 35.939 ;
      RECT 40.975 35.837 43.545 35.893 ;
      RECT 41.021 35.791 43.591 35.847 ;
      RECT 41.067 35.745 43.637 35.801 ;
      RECT 41.113 35.699 43.683 35.755 ;
      RECT 41.159 35.653 43.729 35.709 ;
      RECT 41.205 35.607 43.775 35.663 ;
      RECT 41.251 35.561 43.821 35.617 ;
      RECT 41.297 35.515 43.867 35.571 ;
      RECT 41.343 35.469 43.913 35.525 ;
      RECT 41.389 35.423 43.959 35.479 ;
      RECT 41.435 35.377 44.005 35.433 ;
      RECT 41.481 35.331 44.051 35.387 ;
      RECT 41.527 35.285 44.097 35.341 ;
      RECT 41.573 35.239 44.143 35.295 ;
      RECT 41.619 35.193 44.189 35.249 ;
      RECT 41.665 35.147 44.235 35.203 ;
      RECT 41.711 35.101 44.281 35.157 ;
      RECT 41.757 35.055 44.327 35.111 ;
      RECT 41.803 35.009 44.373 35.065 ;
      RECT 41.849 34.963 44.419 35.019 ;
      RECT 41.895 34.917 44.465 34.973 ;
      RECT 41.941 34.871 44.511 34.927 ;
      RECT 41.987 34.825 44.557 34.881 ;
      RECT 42.033 34.779 44.603 34.835 ;
      RECT 42.079 34.733 44.649 34.789 ;
      RECT 42.125 34.687 44.695 34.743 ;
      RECT 42.171 34.641 44.741 34.697 ;
      RECT 42.217 34.595 44.787 34.651 ;
      RECT 42.263 34.549 44.833 34.605 ;
      RECT 42.309 34.503 44.879 34.559 ;
      RECT 42.355 34.457 44.925 34.513 ;
      RECT 42.401 34.411 44.971 34.467 ;
      RECT 42.447 34.365 45.017 34.421 ;
      RECT 42.493 34.319 45.063 34.375 ;
      RECT 42.539 34.273 45.109 34.329 ;
      RECT 42.585 34.227 45.155 34.283 ;
      RECT 42.631 34.181 45.201 34.237 ;
      RECT 42.677 34.135 45.247 34.191 ;
      RECT 42.723 34.089 45.293 34.145 ;
      RECT 42.769 34.043 45.339 34.099 ;
      RECT 42.815 33.997 45.385 34.053 ;
      RECT 42.861 33.951 45.431 34.007 ;
      RECT 42.907 33.905 45.477 33.961 ;
      RECT 42.953 33.859 45.523 33.915 ;
      RECT 42.999 33.813 45.569 33.869 ;
      RECT 43.045 33.767 45.615 33.823 ;
      RECT 43.091 33.721 45.661 33.777 ;
      RECT 43.137 33.675 45.707 33.731 ;
      RECT 43.183 33.629 45.753 33.685 ;
      RECT 43.229 33.583 45.799 33.639 ;
      RECT 43.275 33.537 45.845 33.593 ;
      RECT 43.321 33.491 45.891 33.547 ;
      RECT 43.367 33.445 45.937 33.501 ;
      RECT 43.413 33.399 45.983 33.455 ;
      RECT 43.459 33.353 46.029 33.409 ;
      RECT 43.505 33.307 46.075 33.363 ;
      RECT 43.551 33.261 46.121 33.317 ;
      RECT 43.597 33.215 46.167 33.271 ;
      RECT 43.643 33.169 46.213 33.225 ;
      RECT 43.689 33.123 46.259 33.179 ;
      RECT 43.735 33.077 46.305 33.133 ;
      RECT 43.781 33.031 46.351 33.087 ;
      RECT 43.827 32.985 46.397 33.041 ;
      RECT 43.873 32.939 46.443 32.995 ;
      RECT 43.919 32.893 46.489 32.949 ;
      RECT 43.965 32.847 46.535 32.903 ;
      RECT 44.011 32.801 46.581 32.857 ;
      RECT 44.057 32.755 46.627 32.811 ;
      RECT 44.103 32.709 46.673 32.765 ;
      RECT 44.149 32.663 46.719 32.719 ;
      RECT 44.195 32.617 46.765 32.673 ;
      RECT 44.241 32.571 46.811 32.627 ;
      RECT 44.287 32.525 46.857 32.581 ;
      RECT 44.333 32.479 46.903 32.535 ;
      RECT 44.379 32.433 46.949 32.489 ;
      RECT 44.425 32.387 46.995 32.443 ;
      RECT 44.471 32.341 47.041 32.397 ;
      RECT 44.517 32.295 47.087 32.351 ;
      RECT 44.563 32.249 47.133 32.305 ;
      RECT 44.609 32.203 47.179 32.259 ;
      RECT 44.655 32.157 47.225 32.213 ;
      RECT 44.701 32.111 47.271 32.167 ;
      RECT 44.747 32.065 47.317 32.121 ;
      RECT 44.793 32.019 47.363 32.075 ;
      RECT 44.839 31.973 47.409 32.029 ;
      RECT 44.885 31.927 47.455 31.983 ;
      RECT 44.931 31.881 47.501 31.937 ;
      RECT 44.977 31.835 47.547 31.891 ;
      RECT 45.023 31.789 47.593 31.845 ;
      RECT 45.069 31.743 47.639 31.799 ;
      RECT 45.115 31.697 47.685 31.753 ;
      RECT 45.161 31.651 47.731 31.707 ;
      RECT 45.207 31.605 47.777 31.661 ;
      RECT 45.253 31.559 47.823 31.615 ;
      RECT 45.299 31.513 47.869 31.569 ;
      RECT 45.345 31.467 47.915 31.523 ;
      RECT 45.391 31.421 47.961 31.477 ;
      RECT 45.437 31.375 48.007 31.431 ;
      RECT 45.483 31.329 48.053 31.385 ;
      RECT 45.529 31.283 48.099 31.339 ;
      RECT 45.575 31.237 48.145 31.293 ;
      RECT 45.621 31.191 48.191 31.247 ;
      RECT 45.667 31.145 48.237 31.201 ;
      RECT 45.713 31.099 48.283 31.155 ;
      RECT 45.759 31.053 48.329 31.109 ;
      RECT 45.805 31.007 48.375 31.063 ;
      RECT 45.851 30.961 48.421 31.017 ;
      RECT 45.897 30.915 48.467 30.971 ;
      RECT 45.943 30.869 48.513 30.925 ;
      RECT 45.989 30.823 48.559 30.879 ;
      RECT 46.035 30.777 48.605 30.833 ;
      RECT 46.081 30.731 48.651 30.787 ;
      RECT 46.127 30.685 48.697 30.741 ;
      RECT 46.173 30.639 48.743 30.695 ;
      RECT 46.219 30.593 48.789 30.649 ;
      RECT 46.265 30.547 48.835 30.603 ;
      RECT 46.311 30.501 48.881 30.557 ;
      RECT 46.357 30.455 48.927 30.511 ;
      RECT 46.403 30.409 48.973 30.465 ;
      RECT 46.449 30.363 49.019 30.419 ;
      RECT 46.495 30.317 49.065 30.373 ;
      RECT 46.541 30.271 49.111 30.327 ;
      RECT 46.587 30.225 49.157 30.281 ;
      RECT 46.633 30.179 49.203 30.235 ;
      RECT 46.679 30.133 49.249 30.189 ;
      RECT 46.725 30.087 49.295 30.143 ;
      RECT 46.771 30.041 49.341 30.097 ;
      RECT 46.817 29.995 49.387 30.051 ;
      RECT 46.863 29.949 49.433 30.005 ;
      RECT 46.909 29.903 49.479 29.959 ;
      RECT 46.955 29.857 49.525 29.913 ;
      RECT 47.001 29.811 49.571 29.867 ;
      RECT 47.047 29.765 49.617 29.821 ;
      RECT 47.093 29.719 49.663 29.775 ;
      RECT 47.139 29.673 49.709 29.729 ;
      RECT 47.185 29.627 49.755 29.683 ;
      RECT 47.231 29.581 49.801 29.637 ;
      RECT 47.277 29.535 49.847 29.591 ;
      RECT 47.323 29.489 49.893 29.545 ;
      RECT 47.369 29.443 49.939 29.499 ;
      RECT 47.415 29.397 49.985 29.453 ;
      RECT 47.461 29.351 50.031 29.407 ;
      RECT 47.507 29.305 50.077 29.361 ;
      RECT 47.553 29.259 50.123 29.315 ;
      RECT 47.599 29.213 50.169 29.269 ;
      RECT 47.645 29.167 50.215 29.223 ;
      RECT 47.691 29.121 50.261 29.177 ;
      RECT 47.737 29.075 50.307 29.131 ;
      RECT 47.783 29.029 50.353 29.085 ;
      RECT 47.829 28.983 50.399 29.039 ;
      RECT 47.875 28.937 50.445 28.993 ;
      RECT 47.921 28.891 50.491 28.947 ;
      RECT 47.967 28.845 50.537 28.901 ;
      RECT 48.013 28.799 50.583 28.855 ;
      RECT 48.059 28.753 50.629 28.809 ;
      RECT 48.105 28.707 50.675 28.763 ;
      RECT 48.151 28.661 50.721 28.717 ;
      RECT 48.197 28.615 50.767 28.671 ;
      RECT 48.243 28.569 50.813 28.625 ;
      RECT 48.289 28.523 50.859 28.579 ;
      RECT 48.335 28.477 50.905 28.533 ;
      RECT 48.381 28.431 50.951 28.487 ;
      RECT 48.427 28.385 50.997 28.441 ;
      RECT 48.473 28.339 51.043 28.395 ;
      RECT 48.519 28.293 51.089 28.349 ;
      RECT 48.565 28.247 51.135 28.303 ;
      RECT 48.611 28.201 51.181 28.257 ;
      RECT 48.657 28.155 51.227 28.211 ;
      RECT 48.703 28.109 51.273 28.165 ;
      RECT 48.749 28.063 51.319 28.119 ;
      RECT 48.795 28.017 51.365 28.073 ;
      RECT 48.841 27.971 51.411 28.027 ;
      RECT 48.887 27.925 51.457 27.981 ;
      RECT 48.933 27.879 51.503 27.935 ;
      RECT 48.979 27.833 51.549 27.889 ;
      RECT 49.025 27.787 51.595 27.843 ;
      RECT 49.071 27.741 51.641 27.797 ;
      RECT 49.117 27.695 51.687 27.751 ;
      RECT 49.163 27.649 51.733 27.705 ;
      RECT 49.209 27.603 51.779 27.659 ;
      RECT 49.255 27.557 51.825 27.613 ;
      RECT 49.301 27.511 51.871 27.567 ;
      RECT 49.347 27.465 51.917 27.521 ;
      RECT 49.393 27.419 51.963 27.475 ;
      RECT 49.439 27.373 52.009 27.429 ;
      RECT 49.485 27.327 52.055 27.383 ;
      RECT 49.531 27.281 52.101 27.337 ;
      RECT 49.577 27.235 52.147 27.291 ;
      RECT 49.623 27.189 52.193 27.245 ;
      RECT 49.669 27.143 52.239 27.199 ;
      RECT 49.715 27.097 52.285 27.153 ;
      RECT 49.761 27.051 52.331 27.107 ;
      RECT 49.807 27.005 52.377 27.061 ;
      RECT 49.853 26.959 52.423 27.015 ;
      RECT 49.899 26.913 52.469 26.969 ;
      RECT 49.945 26.867 52.515 26.923 ;
      RECT 49.991 26.821 52.561 26.877 ;
      RECT 50.037 26.775 52.607 26.831 ;
      RECT 50.083 26.729 52.653 26.785 ;
      RECT 50.129 26.683 52.699 26.739 ;
      RECT 50.175 26.637 52.745 26.693 ;
      RECT 50.221 26.591 52.791 26.647 ;
      RECT 50.267 26.545 52.837 26.601 ;
      RECT 50.313 26.499 52.883 26.555 ;
      RECT 50.359 26.453 52.929 26.509 ;
      RECT 50.405 26.407 52.975 26.463 ;
      RECT 50.451 26.361 53.021 26.417 ;
      RECT 50.497 26.315 53.067 26.371 ;
      RECT 50.543 26.269 53.113 26.325 ;
      RECT 50.589 26.223 53.159 26.279 ;
      RECT 50.635 26.177 53.205 26.233 ;
      RECT 50.681 26.131 53.251 26.187 ;
      RECT 50.727 26.085 53.297 26.141 ;
      RECT 50.773 26.039 53.343 26.095 ;
      RECT 50.819 25.993 53.389 26.049 ;
      RECT 50.865 25.947 53.435 26.003 ;
      RECT 50.911 25.901 53.481 25.957 ;
      RECT 50.957 25.855 53.527 25.911 ;
      RECT 51.003 25.809 53.573 25.865 ;
      RECT 51.049 25.763 53.619 25.819 ;
      RECT 51.095 25.717 53.665 25.773 ;
      RECT 51.141 25.671 53.711 25.727 ;
      RECT 51.187 25.625 53.757 25.681 ;
      RECT 51.233 25.579 53.803 25.635 ;
      RECT 51.279 25.533 53.849 25.589 ;
      RECT 51.325 25.487 53.895 25.543 ;
      RECT 51.371 25.441 53.941 25.497 ;
      RECT 51.417 25.395 53.987 25.451 ;
      RECT 51.463 25.349 54.033 25.405 ;
      RECT 51.509 25.303 54.079 25.359 ;
      RECT 51.555 25.257 54.125 25.313 ;
      RECT 51.601 25.211 54.171 25.267 ;
      RECT 51.647 25.165 54.217 25.221 ;
      RECT 51.693 25.119 54.263 25.175 ;
      RECT 51.739 25.073 54.309 25.129 ;
      RECT 51.785 25.027 54.355 25.083 ;
      RECT 51.831 24.981 54.401 25.037 ;
      RECT 51.877 24.935 54.447 24.991 ;
      RECT 51.923 24.889 54.493 24.945 ;
      RECT 51.969 24.843 54.539 24.899 ;
      RECT 52.015 24.797 54.585 24.853 ;
      RECT 52.061 24.751 54.631 24.807 ;
      RECT 52.107 24.705 54.677 24.761 ;
      RECT 52.153 24.659 54.723 24.715 ;
      RECT 52.199 24.613 54.769 24.669 ;
      RECT 52.245 24.567 54.815 24.623 ;
      RECT 52.291 24.521 54.861 24.577 ;
      RECT 52.337 24.475 54.907 24.531 ;
      RECT 52.383 24.429 54.953 24.485 ;
      RECT 52.429 24.383 54.999 24.439 ;
      RECT 52.475 24.337 55.045 24.393 ;
      RECT 52.521 24.291 55.091 24.347 ;
      RECT 52.567 24.245 55.137 24.301 ;
      RECT 52.613 24.199 55.183 24.255 ;
      RECT 52.659 24.153 55.229 24.209 ;
      RECT 52.705 24.107 55.275 24.163 ;
      RECT 52.751 24.061 55.321 24.117 ;
      RECT 52.797 24.015 55.367 24.071 ;
      RECT 52.843 23.969 55.413 24.025 ;
      RECT 52.889 23.923 55.459 23.979 ;
      RECT 52.935 23.877 55.505 23.933 ;
      RECT 52.981 23.831 55.551 23.887 ;
      RECT 53.027 23.785 55.597 23.841 ;
      RECT 53.073 23.739 55.643 23.795 ;
      RECT 53.119 23.693 55.689 23.749 ;
      RECT 53.165 23.647 55.735 23.703 ;
      RECT 53.211 23.601 55.781 23.657 ;
      RECT 53.257 23.555 55.827 23.611 ;
      RECT 53.303 23.509 55.873 23.565 ;
      RECT 53.349 23.463 55.919 23.519 ;
      RECT 53.395 23.417 55.965 23.473 ;
      RECT 53.441 23.371 56.011 23.427 ;
      RECT 53.487 23.325 56.057 23.381 ;
      RECT 53.533 23.279 56.103 23.335 ;
      RECT 53.579 23.233 56.149 23.289 ;
      RECT 53.625 23.187 56.195 23.243 ;
      RECT 53.671 23.141 56.241 23.197 ;
      RECT 53.717 23.095 56.287 23.151 ;
      RECT 53.763 23.049 56.333 23.105 ;
      RECT 53.809 23.003 56.379 23.059 ;
      RECT 53.855 22.957 56.425 23.013 ;
      RECT 53.901 22.911 56.471 22.967 ;
      RECT 53.947 22.865 56.517 22.921 ;
      RECT 53.993 22.819 56.563 22.875 ;
      RECT 54.039 22.773 56.609 22.829 ;
      RECT 54.085 22.727 56.655 22.783 ;
      RECT 54.131 22.681 56.701 22.737 ;
      RECT 54.177 22.635 56.747 22.691 ;
      RECT 54.223 22.589 56.793 22.645 ;
      RECT 54.269 22.543 56.839 22.599 ;
      RECT 54.315 22.497 56.885 22.553 ;
      RECT 54.361 22.451 56.931 22.507 ;
      RECT 54.407 22.405 56.977 22.461 ;
      RECT 54.453 22.359 57.023 22.415 ;
      RECT 54.499 22.313 57.069 22.369 ;
      RECT 54.545 22.267 57.115 22.323 ;
      RECT 54.591 22.221 57.161 22.277 ;
      RECT 54.637 22.175 57.207 22.231 ;
      RECT 54.683 22.129 57.253 22.185 ;
      RECT 54.729 22.083 57.299 22.139 ;
      RECT 54.775 22.037 57.345 22.093 ;
      RECT 54.821 21.991 57.391 22.047 ;
      RECT 54.867 21.945 57.437 22.001 ;
      RECT 54.913 21.899 57.483 21.955 ;
      RECT 54.959 21.853 57.529 21.909 ;
      RECT 55.005 21.807 57.575 21.863 ;
      RECT 55.051 21.761 57.621 21.817 ;
      RECT 55.097 21.715 57.667 21.771 ;
      RECT 55.143 21.669 57.713 21.725 ;
      RECT 55.189 21.623 57.759 21.679 ;
      RECT 55.235 21.577 57.805 21.633 ;
      RECT 55.281 21.531 57.851 21.587 ;
      RECT 55.327 21.485 57.897 21.541 ;
      RECT 55.373 21.439 57.943 21.495 ;
      RECT 55.419 21.393 57.989 21.449 ;
      RECT 55.465 21.347 58.035 21.403 ;
      RECT 55.511 21.301 58.081 21.357 ;
      RECT 55.557 21.255 58.127 21.311 ;
      RECT 55.603 21.209 58.173 21.265 ;
      RECT 55.649 21.163 58.219 21.219 ;
      RECT 55.695 21.117 58.265 21.173 ;
      RECT 55.741 21.071 58.311 21.127 ;
      RECT 55.787 21.025 58.357 21.081 ;
      RECT 55.833 20.979 58.403 21.035 ;
      RECT 55.879 20.933 58.449 20.989 ;
      RECT 55.925 20.887 58.495 20.943 ;
      RECT 55.971 20.841 58.541 20.897 ;
      RECT 56.017 20.795 58.587 20.851 ;
      RECT 56.063 20.749 58.633 20.805 ;
      RECT 56.109 20.703 58.679 20.759 ;
      RECT 56.155 20.663 58.725 20.713 ;
      RECT 56.19 20.622 58.771 20.667 ;
      RECT 56.236 20.576 58.817 20.621 ;
      RECT 56.282 20.53 58.863 20.575 ;
      RECT 56.328 20.484 58.909 20.529 ;
      RECT 56.374 20.438 58.955 20.483 ;
      RECT 56.42 20.392 59.001 20.437 ;
      RECT 56.466 20.346 59.047 20.391 ;
      RECT 56.512 20.3 59.093 20.345 ;
      RECT 56.558 20.254 59.139 20.299 ;
      RECT 56.604 20.208 59.185 20.253 ;
      RECT 56.65 20.162 59.231 20.207 ;
      RECT 56.696 20.116 59.277 20.161 ;
      RECT 56.742 20.07 59.323 20.115 ;
      RECT 56.788 20.024 59.369 20.069 ;
      RECT 56.834 19.978 59.415 20.023 ;
      RECT 56.88 19.932 59.461 19.977 ;
      RECT 56.926 19.886 59.507 19.931 ;
      RECT 56.972 19.84 59.553 19.885 ;
      RECT 57.018 19.794 59.599 19.839 ;
      RECT 57.064 19.748 59.645 19.793 ;
      RECT 57.11 19.702 59.691 19.747 ;
      RECT 57.156 19.656 59.737 19.701 ;
      RECT 57.202 19.61 59.783 19.655 ;
      RECT 57.248 19.564 59.829 19.609 ;
      RECT 57.294 19.518 59.875 19.563 ;
      RECT 57.34 19.472 59.921 19.517 ;
      RECT 57.386 19.426 59.967 19.471 ;
      RECT 57.432 19.38 60.013 19.425 ;
      RECT 57.478 19.334 60.059 19.379 ;
      RECT 57.524 19.288 60.105 19.333 ;
      RECT 57.57 19.242 60.151 19.287 ;
      RECT 57.616 19.196 60.197 19.241 ;
      RECT 57.662 19.15 60.243 19.195 ;
      RECT 57.708 19.104 60.289 19.149 ;
      RECT 57.754 19.058 60.335 19.103 ;
      RECT 57.8 19.012 60.381 19.057 ;
      RECT 57.846 18.966 60.427 19.011 ;
      RECT 57.892 18.92 60.473 18.965 ;
      RECT 57.938 18.874 60.519 18.919 ;
      RECT 57.984 18.828 60.565 18.873 ;
      RECT 58.03 18.782 60.611 18.827 ;
      RECT 58.076 18.736 60.657 18.781 ;
      RECT 58.122 18.69 60.703 18.735 ;
      RECT 58.168 18.644 60.749 18.689 ;
      RECT 58.214 18.598 60.795 18.643 ;
      RECT 58.26 18.552 60.841 18.597 ;
      RECT 58.306 18.506 60.887 18.551 ;
      RECT 58.352 18.46 60.933 18.505 ;
      RECT 58.398 18.414 60.979 18.459 ;
      RECT 58.444 18.368 61.025 18.413 ;
      RECT 58.49 18.322 61.071 18.367 ;
      RECT 58.536 18.276 61.117 18.321 ;
      RECT 58.582 18.23 61.163 18.275 ;
      RECT 58.628 18.184 61.209 18.229 ;
      RECT 58.674 18.138 61.255 18.183 ;
      RECT 58.72 18.092 61.301 18.137 ;
      RECT 58.766 18.046 61.347 18.091 ;
      RECT 58.812 18 61.393 18.045 ;
      RECT 58.858 17.954 61.439 17.999 ;
      RECT 58.904 17.908 61.485 17.953 ;
      RECT 58.95 17.862 61.531 17.907 ;
      RECT 58.996 17.816 61.577 17.861 ;
      RECT 59.042 17.77 61.623 17.815 ;
      RECT 59.088 17.724 61.669 17.769 ;
      RECT 59.134 17.678 61.715 17.723 ;
      RECT 59.18 17.632 61.761 17.677 ;
      RECT 59.226 17.586 61.807 17.631 ;
      RECT 59.272 17.54 61.853 17.585 ;
      RECT 59.318 17.494 61.899 17.539 ;
      RECT 59.364 17.448 61.945 17.493 ;
      RECT 59.41 17.402 61.991 17.447 ;
      RECT 59.456 17.356 62.037 17.401 ;
      RECT 59.502 17.31 62.083 17.355 ;
      RECT 59.548 17.264 62.129 17.309 ;
      RECT 59.594 17.218 62.175 17.263 ;
      RECT 59.64 17.172 62.221 17.217 ;
      RECT 59.686 17.126 62.267 17.171 ;
      RECT 59.732 17.08 62.313 17.125 ;
      RECT 59.778 17.034 62.359 17.079 ;
      RECT 59.824 16.988 62.405 17.033 ;
      RECT 59.87 16.942 62.451 16.987 ;
      RECT 59.916 16.896 62.497 16.941 ;
      RECT 59.962 16.85 62.543 16.895 ;
      RECT 60.008 16.804 62.589 16.849 ;
      RECT 61.158 15.675 110 16.825 ;
      RECT 60.054 16.758 110 16.825 ;
      RECT 61.112 15.699 61.163 18.275 ;
      RECT 60.1 16.712 110 16.825 ;
      RECT 61.066 15.746 61.117 18.321 ;
      RECT 60.146 16.666 110 16.825 ;
      RECT 61.02 15.792 61.071 18.367 ;
      RECT 60.192 16.62 110 16.825 ;
      RECT 60.974 15.838 61.025 18.413 ;
      RECT 60.238 16.574 110 16.825 ;
      RECT 60.928 15.884 60.979 18.459 ;
      RECT 60.284 16.528 110 16.825 ;
      RECT 60.882 15.93 60.933 18.505 ;
      RECT 60.33 16.482 110 16.825 ;
      RECT 60.836 15.976 60.887 18.551 ;
      RECT 60.376 16.436 110 16.825 ;
      RECT 60.79 16.022 60.841 18.597 ;
      RECT 60.422 16.39 110 16.825 ;
      RECT 60.744 16.068 60.795 18.643 ;
      RECT 60.468 16.344 110 16.825 ;
      RECT 60.698 16.114 60.749 18.689 ;
      RECT 60.514 16.298 110 16.825 ;
      RECT 60.652 16.16 60.703 18.735 ;
      RECT 60.56 16.252 110 16.825 ;
      RECT 60.606 16.206 60.657 18.781 ;
      RECT 29.175 67.887 30.325 110 ;
      RECT 29.175 67.887 30.371 69.317 ;
      RECT 29.175 67.887 30.417 69.271 ;
      RECT 29.175 67.887 30.463 69.225 ;
      RECT 29.175 67.887 30.509 69.179 ;
      RECT 29.175 67.887 30.555 69.133 ;
      RECT 29.175 67.887 30.601 69.087 ;
      RECT 29.175 67.887 30.647 69.041 ;
      RECT 29.175 67.887 30.693 68.995 ;
      RECT 29.175 67.887 30.739 68.949 ;
      RECT 29.175 67.887 30.785 68.903 ;
      RECT 29.175 67.887 30.831 68.857 ;
      RECT 29.175 67.887 30.877 68.811 ;
      RECT 29.175 67.887 30.923 68.765 ;
      RECT 29.175 67.887 30.969 68.719 ;
      RECT 29.175 67.887 31.015 68.673 ;
      RECT 29.175 67.887 31.061 68.627 ;
      RECT 29.175 67.887 31.107 68.581 ;
      RECT 29.175 67.887 31.153 68.535 ;
      RECT 29.175 67.887 31.199 68.489 ;
      RECT 29.175 67.887 31.245 68.443 ;
      RECT 29.175 67.887 31.291 68.397 ;
      RECT 29.175 67.887 31.337 68.351 ;
      RECT 29.175 67.887 31.383 68.305 ;
      RECT 29.175 67.887 31.429 68.259 ;
      RECT 29.175 67.887 31.475 68.213 ;
      RECT 29.175 67.887 31.521 68.167 ;
      RECT 29.175 67.887 31.567 68.121 ;
      RECT 29.175 67.887 31.613 68.075 ;
      RECT 29.175 67.887 31.659 68.029 ;
      RECT 29.175 67.887 31.705 67.983 ;
      RECT 29.175 67.887 31.751 67.937 ;
      RECT 29.221 67.841 31.797 67.891 ;
      RECT 29.267 67.795 31.843 67.845 ;
      RECT 29.313 67.749 31.889 67.799 ;
      RECT 29.359 67.703 31.935 67.753 ;
      RECT 29.405 67.657 31.981 67.707 ;
      RECT 29.451 67.611 32.027 67.661 ;
      RECT 29.497 67.565 32.073 67.615 ;
      RECT 29.543 67.519 32.119 67.569 ;
      RECT 29.589 67.473 32.165 67.523 ;
      RECT 29.635 67.427 32.211 67.477 ;
      RECT 29.681 67.381 32.257 67.431 ;
      RECT 29.727 67.335 32.303 67.385 ;
      RECT 29.773 67.289 32.349 67.339 ;
      RECT 29.819 67.243 32.395 67.293 ;
      RECT 29.865 67.197 32.441 67.247 ;
      RECT 29.911 67.151 32.487 67.201 ;
      RECT 29.957 67.105 32.533 67.155 ;
      RECT 30.003 67.059 32.579 67.109 ;
      RECT 30.049 67.013 32.625 67.063 ;
      RECT 30.095 66.967 32.671 67.017 ;
      RECT 30.141 66.921 32.717 66.971 ;
      RECT 30.187 66.875 32.763 66.925 ;
      RECT 30.233 66.829 32.809 66.879 ;
      RECT 30.279 66.783 32.855 66.833 ;
      RECT 30.325 66.737 32.901 66.787 ;
      RECT 30.371 66.691 32.947 66.741 ;
      RECT 30.417 66.645 32.993 66.695 ;
      RECT 30.463 66.599 33.039 66.649 ;
      RECT 30.509 66.553 33.085 66.603 ;
      RECT 30.555 66.507 33.131 66.557 ;
      RECT 30.601 66.461 33.177 66.511 ;
      RECT 30.647 66.415 33.223 66.465 ;
      RECT 30.693 66.369 33.269 66.419 ;
      RECT 30.739 66.323 33.315 66.373 ;
      RECT 30.785 66.277 33.361 66.327 ;
      RECT 30.831 66.231 33.407 66.281 ;
      RECT 30.877 66.185 33.453 66.235 ;
      RECT 30.923 66.139 33.499 66.189 ;
      RECT 30.969 66.093 33.545 66.143 ;
      RECT 31.015 66.047 33.591 66.097 ;
      RECT 31.061 66.001 33.637 66.051 ;
      RECT 31.107 65.955 33.683 66.005 ;
      RECT 31.153 65.909 33.729 65.959 ;
      RECT 31.199 65.863 33.775 65.913 ;
      RECT 31.245 65.817 33.821 65.867 ;
      RECT 31.291 65.771 33.867 65.821 ;
      RECT 31.337 65.725 33.913 65.775 ;
      RECT 31.383 65.679 33.959 65.729 ;
      RECT 31.429 65.633 34.005 65.683 ;
      RECT 31.475 65.587 34.051 65.637 ;
      RECT 31.521 65.541 34.097 65.591 ;
      RECT 31.567 65.495 34.143 65.545 ;
      RECT 31.613 65.449 34.189 65.499 ;
      RECT 31.659 65.403 34.235 65.453 ;
      RECT 31.705 65.357 34.281 65.407 ;
      RECT 31.751 65.311 34.327 65.361 ;
      RECT 31.797 65.265 34.373 65.315 ;
      RECT 31.843 65.219 34.419 65.269 ;
      RECT 31.889 65.173 34.465 65.223 ;
      RECT 31.935 65.127 34.511 65.177 ;
      RECT 31.981 65.081 34.557 65.131 ;
      RECT 32.027 65.035 34.603 65.085 ;
      RECT 32.073 64.989 34.649 65.039 ;
      RECT 32.119 64.943 34.695 64.993 ;
      RECT 32.165 64.897 34.741 64.947 ;
      RECT 32.211 64.851 34.787 64.901 ;
      RECT 32.257 64.805 34.833 64.855 ;
      RECT 32.303 64.759 34.879 64.809 ;
      RECT 32.349 64.713 34.925 64.763 ;
      RECT 32.395 64.667 34.971 64.717 ;
      RECT 32.441 64.621 35.017 64.671 ;
      RECT 32.487 64.575 35.063 64.625 ;
      RECT 32.533 64.529 35.109 64.579 ;
      RECT 32.579 64.483 35.155 64.533 ;
      RECT 32.625 64.437 35.201 64.487 ;
      RECT 32.671 64.391 35.247 64.441 ;
      RECT 32.717 64.345 35.293 64.395 ;
      RECT 32.763 64.299 35.339 64.349 ;
      RECT 32.809 64.253 35.385 64.303 ;
      RECT 32.855 64.207 35.431 64.257 ;
      RECT 32.901 64.161 35.477 64.211 ;
      RECT 32.947 64.115 35.523 64.165 ;
      RECT 32.993 64.069 35.569 64.119 ;
      RECT 33.039 64.023 35.615 64.073 ;
      RECT 33.085 63.977 35.661 64.027 ;
      RECT 33.131 63.931 35.707 63.981 ;
      RECT 33.177 63.885 35.753 63.935 ;
      RECT 33.223 63.839 35.799 63.889 ;
      RECT 33.269 63.793 35.845 63.843 ;
      RECT 33.315 63.747 35.891 63.797 ;
      RECT 33.361 63.701 35.937 63.751 ;
      RECT 33.407 63.655 35.983 63.705 ;
      RECT 33.453 63.609 36.029 63.659 ;
      RECT 33.499 63.563 36.075 63.613 ;
      RECT 33.545 63.517 36.121 63.567 ;
      RECT 33.591 63.471 36.167 63.521 ;
      RECT 33.637 63.425 36.213 63.475 ;
      RECT 33.683 63.379 36.259 63.429 ;
      RECT 33.729 63.333 36.305 63.383 ;
      RECT 33.775 63.287 36.351 63.337 ;
      RECT 33.821 63.241 36.397 63.291 ;
      RECT 33.867 63.195 36.443 63.245 ;
      RECT 33.913 63.149 36.489 63.199 ;
      RECT 33.959 63.103 36.535 63.153 ;
      RECT 34.005 63.057 36.581 63.107 ;
      RECT 34.051 63.011 36.627 63.061 ;
      RECT 34.097 62.965 36.673 63.015 ;
      RECT 34.143 62.919 36.719 62.969 ;
      RECT 34.189 62.873 36.765 62.923 ;
      RECT 34.235 62.827 36.811 62.877 ;
      RECT 34.281 62.781 36.857 62.831 ;
      RECT 34.327 62.735 36.903 62.785 ;
      RECT 34.373 62.689 36.949 62.739 ;
      RECT 34.419 62.643 36.995 62.693 ;
      RECT 34.465 62.597 37.041 62.647 ;
      RECT 34.511 62.551 37.087 62.601 ;
      RECT 34.557 62.505 37.133 62.555 ;
      RECT 34.603 62.459 37.179 62.509 ;
      RECT 34.649 62.413 37.225 62.463 ;
      RECT 34.695 62.367 37.271 62.417 ;
      RECT 34.741 62.321 37.317 62.371 ;
      RECT 34.787 62.275 37.363 62.325 ;
      RECT 34.833 62.229 37.409 62.279 ;
      RECT 34.879 62.183 37.455 62.233 ;
      RECT 34.925 62.137 37.501 62.187 ;
      RECT 34.971 62.091 37.547 62.141 ;
      RECT 35.017 62.045 37.593 62.095 ;
      RECT 35.063 61.999 37.639 62.049 ;
      RECT 35.109 61.953 37.685 62.003 ;
      RECT 35.155 61.907 37.731 61.957 ;
      RECT 35.201 61.861 37.777 61.911 ;
      RECT 35.247 61.815 37.823 61.865 ;
      RECT 35.293 61.769 37.869 61.819 ;
      RECT 35.339 61.723 37.915 61.773 ;
      RECT 35.385 61.677 37.961 61.727 ;
      RECT 35.431 61.631 38.007 61.681 ;
      RECT 35.477 61.585 38.053 61.635 ;
      RECT 35.523 61.539 38.099 61.589 ;
      RECT 35.569 61.493 38.145 61.543 ;
      RECT 35.615 61.447 38.191 61.497 ;
      RECT 35.661 61.401 38.237 61.451 ;
      RECT 35.707 61.355 38.283 61.405 ;
      RECT 35.753 61.309 38.329 61.359 ;
      RECT 35.799 61.263 38.375 61.313 ;
      RECT 35.845 61.217 38.421 61.267 ;
      RECT 35.891 61.171 38.467 61.221 ;
      RECT 35.937 61.125 38.513 61.175 ;
      RECT 35.983 61.079 38.559 61.129 ;
      RECT 36.029 61.033 38.605 61.083 ;
      RECT 36.075 60.987 38.651 61.037 ;
      RECT 36.121 60.941 38.697 60.991 ;
      RECT 36.167 60.895 38.743 60.945 ;
      RECT 36.213 60.849 38.789 60.899 ;
      RECT 36.259 60.803 38.835 60.853 ;
      RECT 36.305 60.757 38.881 60.807 ;
      RECT 36.351 60.711 38.927 60.761 ;
      RECT 36.397 60.665 38.973 60.715 ;
      RECT 36.443 60.619 39.019 60.669 ;
      RECT 36.489 60.573 39.065 60.623 ;
      RECT 36.535 60.527 39.111 60.577 ;
      RECT 36.581 60.481 39.157 60.531 ;
      RECT 36.627 60.435 39.203 60.485 ;
      RECT 36.673 60.389 39.249 60.439 ;
      RECT 36.719 60.343 39.295 60.393 ;
      RECT 36.765 60.297 39.341 60.347 ;
      RECT 36.811 60.251 39.387 60.301 ;
      RECT 36.857 60.205 39.433 60.255 ;
      RECT 36.903 60.159 39.479 60.209 ;
      RECT 36.949 60.113 39.525 60.163 ;
      RECT 36.995 60.067 39.571 60.117 ;
      RECT 37.041 60.021 39.617 60.071 ;
      RECT 37.087 59.975 39.663 60.025 ;
      RECT 37.133 59.929 39.709 59.979 ;
      RECT 37.179 59.883 39.755 59.933 ;
      RECT 37.225 59.837 39.801 59.887 ;
      RECT 37.271 59.791 39.847 59.841 ;
      RECT 37.317 59.745 39.893 59.795 ;
      RECT 37.363 59.699 39.939 59.749 ;
      RECT 37.409 59.653 39.985 59.703 ;
      RECT 37.455 59.607 40.031 59.657 ;
      RECT 37.501 59.561 40.077 59.611 ;
      RECT 37.547 59.515 40.123 59.565 ;
      RECT 37.593 59.469 40.169 59.519 ;
      RECT 37.639 59.423 40.215 59.473 ;
      RECT 37.685 59.377 40.261 59.427 ;
      RECT 37.731 59.331 40.307 59.381 ;
      RECT 37.777 59.285 40.353 59.335 ;
      RECT 37.823 59.239 40.399 59.289 ;
      RECT 37.869 59.193 40.445 59.243 ;
      RECT 37.915 59.147 40.491 59.197 ;
      RECT 37.961 59.101 40.537 59.151 ;
      RECT 38.007 59.055 40.583 59.105 ;
      RECT 38.053 59.009 40.629 59.059 ;
      RECT 38.099 58.963 40.675 59.013 ;
      RECT 38.145 58.917 40.721 58.967 ;
      RECT 38.191 58.871 40.767 58.921 ;
      RECT 38.237 58.825 40.813 58.875 ;
      RECT 38.283 58.779 40.859 58.829 ;
      RECT 38.329 58.733 40.905 58.783 ;
      RECT 38.375 58.687 40.951 58.737 ;
      RECT 38.421 58.641 40.997 58.691 ;
      RECT 38.467 58.595 41.043 58.645 ;
      RECT 38.513 58.549 41.089 58.599 ;
      RECT 38.559 58.503 41.135 58.553 ;
      RECT 38.605 58.457 41.181 58.507 ;
      RECT 38.651 58.411 41.227 58.461 ;
      RECT 38.697 58.365 41.273 58.415 ;
      RECT 38.743 58.319 41.319 58.369 ;
      RECT 38.789 58.273 41.365 58.323 ;
      RECT 38.835 58.227 41.411 58.277 ;
      RECT 38.881 58.181 41.457 58.231 ;
      RECT 38.927 58.135 41.503 58.185 ;
      RECT 38.973 58.089 41.549 58.139 ;
      RECT 39.019 58.043 41.595 58.093 ;
      RECT 39.065 57.997 41.641 58.047 ;
      RECT 39.111 57.951 41.687 58.001 ;
      RECT 39.157 57.905 41.733 57.955 ;
      RECT 39.203 57.859 41.779 57.909 ;
      RECT 39.249 57.813 41.825 57.863 ;
      RECT 39.295 57.767 41.871 57.817 ;
      RECT 39.341 57.721 41.917 57.771 ;
      RECT 39.387 57.675 41.963 57.725 ;
      RECT 39.433 57.629 42.009 57.679 ;
      RECT 39.479 57.583 42.055 57.633 ;
      RECT 39.525 57.537 42.101 57.587 ;
      RECT 39.571 57.491 42.147 57.541 ;
      RECT 39.617 57.445 42.193 57.495 ;
      RECT 39.663 57.399 42.239 57.449 ;
      RECT 39.709 57.353 42.285 57.403 ;
      RECT 39.755 57.307 42.325 57.36 ;
      RECT 39.801 57.261 42.371 57.317 ;
      RECT 39.847 57.215 42.417 57.271 ;
      RECT 39.893 57.169 42.463 57.225 ;
      RECT 39.939 57.123 42.509 57.179 ;
      RECT 39.985 57.077 42.555 57.133 ;
      RECT 40.031 57.031 42.601 57.087 ;
      RECT 40.077 56.985 42.647 57.041 ;
      RECT 40.123 56.939 42.693 56.995 ;
      RECT 40.169 56.893 42.739 56.949 ;
      RECT 40.215 56.847 42.785 56.903 ;
      RECT 40.261 56.801 42.831 56.857 ;
      RECT 40.307 56.755 42.877 56.811 ;
      RECT 40.353 56.709 42.923 56.765 ;
      RECT 40.399 56.663 42.969 56.719 ;
      RECT 40.445 56.617 43.015 56.673 ;
      RECT 40.491 56.571 43.061 56.627 ;
      RECT 40.537 56.525 43.107 56.581 ;
      RECT 40.583 56.479 43.153 56.535 ;
      RECT 40.629 56.433 43.199 56.489 ;
      RECT 40.675 56.387 43.245 56.443 ;
      RECT 40.721 56.341 43.291 56.397 ;
      RECT 40.767 56.295 43.337 56.351 ;
      RECT 40.813 56.249 43.383 56.305 ;
      RECT 40.859 56.203 43.429 56.259 ;
      RECT 40.905 56.157 43.475 56.213 ;
      RECT 40.951 56.111 43.521 56.167 ;
      RECT 40.997 56.065 43.567 56.121 ;
      RECT 41.043 56.019 43.613 56.075 ;
      RECT 41.089 55.973 43.659 56.029 ;
      RECT 41.135 55.927 43.705 55.983 ;
      RECT 41.181 55.881 43.751 55.937 ;
      RECT 41.227 55.835 43.797 55.891 ;
      RECT 41.273 55.789 43.843 55.845 ;
      RECT 41.319 55.743 43.889 55.799 ;
      RECT 41.365 55.697 43.935 55.753 ;
      RECT 41.411 55.651 43.981 55.707 ;
      RECT 41.457 55.605 44.027 55.661 ;
      RECT 41.503 55.559 44.073 55.615 ;
      RECT 41.549 55.513 44.119 55.569 ;
      RECT 41.595 55.467 44.165 55.523 ;
      RECT 41.641 55.421 44.211 55.477 ;
      RECT 41.687 55.375 44.257 55.431 ;
      RECT 41.733 55.329 44.303 55.385 ;
      RECT 41.779 55.283 44.349 55.339 ;
      RECT 41.825 55.237 44.395 55.293 ;
      RECT 41.871 55.191 44.441 55.247 ;
      RECT 41.917 55.145 44.487 55.201 ;
      RECT 41.963 55.099 44.533 55.155 ;
      RECT 42.009 55.053 44.579 55.109 ;
      RECT 42.055 55.007 44.625 55.063 ;
      RECT 42.101 54.961 44.671 55.017 ;
      RECT 42.147 54.915 44.717 54.971 ;
      RECT 42.193 54.869 44.763 54.925 ;
      RECT 42.239 54.823 44.809 54.879 ;
      RECT 42.285 54.777 44.855 54.833 ;
      RECT 42.331 54.731 44.901 54.787 ;
      RECT 42.377 54.685 44.947 54.741 ;
      RECT 42.423 54.639 44.993 54.695 ;
      RECT 42.469 54.593 45.039 54.649 ;
      RECT 42.515 54.547 45.085 54.603 ;
      RECT 42.561 54.501 45.131 54.557 ;
      RECT 42.607 54.455 45.177 54.511 ;
      RECT 42.653 54.409 45.223 54.465 ;
      RECT 42.699 54.363 45.269 54.419 ;
      RECT 42.745 54.317 45.315 54.373 ;
      RECT 42.791 54.271 45.361 54.327 ;
      RECT 42.837 54.225 45.407 54.281 ;
      RECT 42.883 54.179 45.453 54.235 ;
      RECT 42.929 54.133 45.499 54.189 ;
      RECT 42.975 54.087 45.545 54.143 ;
      RECT 43.021 54.041 45.591 54.097 ;
      RECT 43.067 53.995 45.637 54.051 ;
      RECT 43.113 53.949 45.683 54.005 ;
      RECT 43.159 53.903 45.729 53.959 ;
      RECT 43.205 53.857 45.775 53.913 ;
      RECT 43.251 53.811 45.821 53.867 ;
      RECT 43.297 53.765 45.867 53.821 ;
      RECT 43.343 53.719 45.913 53.775 ;
      RECT 43.389 53.673 45.959 53.729 ;
      RECT 43.435 53.627 46.005 53.683 ;
      RECT 43.481 53.581 46.051 53.637 ;
      RECT 43.527 53.535 46.097 53.591 ;
      RECT 43.573 53.489 46.143 53.545 ;
      RECT 43.619 53.443 46.189 53.499 ;
      RECT 43.665 53.397 46.235 53.453 ;
      RECT 43.711 53.351 46.281 53.407 ;
      RECT 43.757 53.305 46.327 53.361 ;
      RECT 43.803 53.259 46.373 53.315 ;
      RECT 43.849 53.213 46.419 53.269 ;
      RECT 43.895 53.167 46.465 53.223 ;
      RECT 43.941 53.121 46.511 53.177 ;
      RECT 43.987 53.075 46.557 53.131 ;
      RECT 44.033 53.029 46.603 53.085 ;
      RECT 44.079 52.983 46.649 53.039 ;
      RECT 44.125 52.937 46.695 52.993 ;
      RECT 44.171 52.891 46.741 52.947 ;
      RECT 44.217 52.845 46.787 52.901 ;
      RECT 44.263 52.799 46.833 52.855 ;
      RECT 44.309 52.753 46.879 52.809 ;
      RECT 44.355 52.707 46.925 52.763 ;
      RECT 44.401 52.661 46.971 52.717 ;
      RECT 44.447 52.615 47.017 52.671 ;
      RECT 44.493 52.569 47.063 52.625 ;
      RECT 44.539 52.523 47.109 52.579 ;
      RECT 44.585 52.477 47.155 52.533 ;
      RECT 44.631 52.431 47.201 52.487 ;
      RECT 44.677 52.385 47.247 52.441 ;
      RECT 44.723 52.339 47.293 52.395 ;
      RECT 44.769 52.293 47.339 52.349 ;
      RECT 44.815 52.247 47.385 52.303 ;
      RECT 44.861 52.201 47.431 52.257 ;
      RECT 44.907 52.155 47.477 52.211 ;
      RECT 44.953 52.109 47.523 52.165 ;
      RECT 44.999 52.063 47.569 52.119 ;
      RECT 45.045 52.017 47.615 52.073 ;
      RECT 45.091 51.971 47.661 52.027 ;
      RECT 45.137 51.925 47.707 51.981 ;
      RECT 45.183 51.879 47.753 51.935 ;
      RECT 45.229 51.833 47.799 51.889 ;
      RECT 45.275 51.787 47.845 51.843 ;
      RECT 45.321 51.741 47.891 51.797 ;
      RECT 45.367 51.695 47.937 51.751 ;
      RECT 45.413 51.649 47.983 51.705 ;
      RECT 45.459 51.603 48.029 51.659 ;
      RECT 45.505 51.557 48.075 51.613 ;
      RECT 45.551 51.511 48.121 51.567 ;
      RECT 45.597 51.465 48.167 51.521 ;
      RECT 45.643 51.419 48.213 51.475 ;
      RECT 45.689 51.373 48.259 51.429 ;
      RECT 45.735 51.327 48.305 51.383 ;
      RECT 45.781 51.281 48.351 51.337 ;
      RECT 45.827 51.235 48.397 51.291 ;
      RECT 45.873 51.189 48.443 51.245 ;
      RECT 45.919 51.143 48.489 51.199 ;
      RECT 45.965 51.097 48.535 51.153 ;
      RECT 46.011 51.051 48.581 51.107 ;
      RECT 46.057 51.005 48.627 51.061 ;
      RECT 46.103 50.959 48.673 51.015 ;
      RECT 46.149 50.913 48.719 50.969 ;
      RECT 46.195 50.867 48.765 50.923 ;
      RECT 46.241 50.821 48.811 50.877 ;
      RECT 46.287 50.775 48.857 50.831 ;
      RECT 46.333 50.729 48.903 50.785 ;
      RECT 46.379 50.683 48.949 50.739 ;
      RECT 46.425 50.637 48.995 50.693 ;
      RECT 46.471 50.591 49.041 50.647 ;
      RECT 46.517 50.545 49.087 50.601 ;
      RECT 46.563 50.499 49.133 50.555 ;
      RECT 46.609 50.453 49.179 50.509 ;
      RECT 46.655 50.407 49.225 50.463 ;
      RECT 46.701 50.361 49.271 50.417 ;
      RECT 46.747 50.315 49.317 50.371 ;
      RECT 46.793 50.269 49.363 50.325 ;
      RECT 46.839 50.223 49.409 50.279 ;
      RECT 46.885 50.177 49.455 50.233 ;
      RECT 46.931 50.131 49.501 50.187 ;
      RECT 46.977 50.085 49.547 50.141 ;
      RECT 47.023 50.039 49.593 50.095 ;
      RECT 47.069 49.993 49.639 50.049 ;
      RECT 47.115 49.947 49.685 50.003 ;
      RECT 47.161 49.901 49.731 49.957 ;
      RECT 47.207 49.855 49.777 49.911 ;
      RECT 47.253 49.809 49.823 49.865 ;
      RECT 47.299 49.763 49.869 49.819 ;
      RECT 47.345 49.717 49.915 49.773 ;
      RECT 47.391 49.671 49.961 49.727 ;
      RECT 47.437 49.625 50.007 49.681 ;
      RECT 47.483 49.579 50.053 49.635 ;
      RECT 47.529 49.533 50.099 49.589 ;
      RECT 47.575 49.487 50.145 49.543 ;
      RECT 47.621 49.441 50.191 49.497 ;
      RECT 47.667 49.395 50.237 49.451 ;
      RECT 47.713 49.349 50.283 49.405 ;
      RECT 47.759 49.303 50.329 49.359 ;
      RECT 47.805 49.257 50.375 49.313 ;
      RECT 47.851 49.211 50.421 49.267 ;
      RECT 47.897 49.165 50.467 49.221 ;
      RECT 47.943 49.119 50.513 49.175 ;
      RECT 47.989 49.073 50.559 49.129 ;
      RECT 48.035 49.027 50.605 49.083 ;
      RECT 48.081 48.981 50.651 49.037 ;
      RECT 48.127 48.935 50.697 48.991 ;
      RECT 48.173 48.889 50.743 48.945 ;
      RECT 48.219 48.843 50.789 48.899 ;
      RECT 48.265 48.797 50.835 48.853 ;
      RECT 48.311 48.751 50.881 48.807 ;
      RECT 48.357 48.705 50.927 48.761 ;
      RECT 48.403 48.659 50.973 48.715 ;
      RECT 48.449 48.613 51.019 48.669 ;
      RECT 48.495 48.567 51.065 48.623 ;
      RECT 48.541 48.521 51.111 48.577 ;
      RECT 48.587 48.475 51.157 48.531 ;
      RECT 48.633 48.429 51.203 48.485 ;
      RECT 48.679 48.383 51.249 48.439 ;
      RECT 48.725 48.337 51.295 48.393 ;
      RECT 48.771 48.291 51.341 48.347 ;
      RECT 48.817 48.245 51.387 48.301 ;
      RECT 48.863 48.199 51.433 48.255 ;
      RECT 48.909 48.153 51.479 48.209 ;
      RECT 48.955 48.107 51.525 48.163 ;
      RECT 49.001 48.061 51.571 48.117 ;
      RECT 49.047 48.015 51.617 48.071 ;
      RECT 49.093 47.969 51.663 48.025 ;
      RECT 49.139 47.923 51.709 47.979 ;
      RECT 49.185 47.877 51.755 47.933 ;
      RECT 49.231 47.831 51.801 47.887 ;
      RECT 49.277 47.785 51.847 47.841 ;
      RECT 49.323 47.739 51.893 47.795 ;
      RECT 49.369 47.693 51.939 47.749 ;
      RECT 49.415 47.647 51.985 47.703 ;
      RECT 49.461 47.601 52.031 47.657 ;
      RECT 49.507 47.555 52.077 47.611 ;
      RECT 49.553 47.509 52.123 47.565 ;
      RECT 49.599 47.463 52.169 47.519 ;
      RECT 49.645 47.417 52.215 47.473 ;
      RECT 49.691 47.371 52.261 47.427 ;
      RECT 49.737 47.325 52.307 47.381 ;
      RECT 49.783 47.279 52.353 47.335 ;
      RECT 49.829 47.233 52.399 47.289 ;
      RECT 49.875 47.187 52.445 47.243 ;
      RECT 49.921 47.141 52.491 47.197 ;
      RECT 49.967 47.095 52.537 47.151 ;
      RECT 50.013 47.049 52.583 47.105 ;
      RECT 50.059 47.003 52.629 47.059 ;
      RECT 50.105 46.957 52.675 47.013 ;
      RECT 50.151 46.911 52.721 46.967 ;
      RECT 50.197 46.865 52.767 46.921 ;
      RECT 50.243 46.819 52.813 46.875 ;
      RECT 50.289 46.773 52.859 46.829 ;
      RECT 50.335 46.727 52.905 46.783 ;
      RECT 50.381 46.681 52.951 46.737 ;
      RECT 50.427 46.635 52.997 46.691 ;
      RECT 50.473 46.589 53.043 46.645 ;
      RECT 50.519 46.543 53.089 46.599 ;
      RECT 50.565 46.497 53.135 46.553 ;
      RECT 50.611 46.451 53.181 46.507 ;
      RECT 50.657 46.405 53.227 46.461 ;
      RECT 50.703 46.359 53.273 46.415 ;
      RECT 50.749 46.313 53.319 46.369 ;
      RECT 50.795 46.267 53.365 46.323 ;
      RECT 50.841 46.221 53.411 46.277 ;
      RECT 50.887 46.175 53.457 46.231 ;
      RECT 50.933 46.129 53.503 46.185 ;
      RECT 50.979 46.083 53.549 46.139 ;
      RECT 51.025 46.037 53.595 46.093 ;
      RECT 51.071 45.991 53.641 46.047 ;
      RECT 51.117 45.945 53.687 46.001 ;
      RECT 51.163 45.899 53.733 45.955 ;
      RECT 51.209 45.853 53.779 45.909 ;
      RECT 51.255 45.807 53.825 45.863 ;
      RECT 51.301 45.761 53.871 45.817 ;
      RECT 51.347 45.715 53.917 45.771 ;
      RECT 51.393 45.669 53.963 45.725 ;
      RECT 51.439 45.623 54.009 45.679 ;
      RECT 51.485 45.577 54.055 45.633 ;
      RECT 51.531 45.531 54.101 45.587 ;
      RECT 51.577 45.485 54.147 45.541 ;
      RECT 51.623 45.439 54.193 45.495 ;
      RECT 51.669 45.393 54.239 45.449 ;
      RECT 51.715 45.347 54.285 45.403 ;
      RECT 51.761 45.301 54.331 45.357 ;
      RECT 51.807 45.255 54.377 45.311 ;
      RECT 51.853 45.209 54.423 45.265 ;
      RECT 51.899 45.163 54.469 45.219 ;
      RECT 51.945 45.117 54.515 45.173 ;
      RECT 51.991 45.071 54.561 45.127 ;
      RECT 52.037 45.025 54.607 45.081 ;
      RECT 52.083 44.979 54.653 45.035 ;
      RECT 52.129 44.933 54.699 44.989 ;
      RECT 52.175 44.887 54.745 44.943 ;
      RECT 52.221 44.841 54.791 44.897 ;
      RECT 52.267 44.795 54.837 44.851 ;
      RECT 52.313 44.749 54.883 44.805 ;
      RECT 52.359 44.703 54.929 44.759 ;
      RECT 52.405 44.657 54.975 44.713 ;
      RECT 52.451 44.611 55.021 44.667 ;
      RECT 52.497 44.565 55.067 44.621 ;
      RECT 52.543 44.519 55.113 44.575 ;
      RECT 52.589 44.473 55.159 44.529 ;
      RECT 52.635 44.427 55.205 44.483 ;
      RECT 52.681 44.381 55.251 44.437 ;
      RECT 52.727 44.335 55.297 44.391 ;
      RECT 52.773 44.289 55.343 44.345 ;
      RECT 52.819 44.243 55.389 44.299 ;
      RECT 52.865 44.197 55.435 44.253 ;
      RECT 52.911 44.151 55.481 44.207 ;
      RECT 52.957 44.105 55.527 44.161 ;
      RECT 53.003 44.059 55.573 44.115 ;
      RECT 53.049 44.013 55.619 44.069 ;
      RECT 53.095 43.967 55.665 44.023 ;
      RECT 53.141 43.921 55.711 43.977 ;
      RECT 53.187 43.875 55.757 43.931 ;
      RECT 53.233 43.829 55.803 43.885 ;
      RECT 53.279 43.783 55.849 43.839 ;
      RECT 53.325 43.737 55.895 43.793 ;
      RECT 53.371 43.691 55.941 43.747 ;
      RECT 53.417 43.645 55.987 43.701 ;
      RECT 53.463 43.599 56.033 43.655 ;
      RECT 53.509 43.553 56.079 43.609 ;
      RECT 53.555 43.507 56.125 43.563 ;
      RECT 53.601 43.461 56.171 43.517 ;
      RECT 53.647 43.415 56.217 43.471 ;
      RECT 53.693 43.369 56.263 43.425 ;
      RECT 53.739 43.323 56.309 43.379 ;
      RECT 53.785 43.277 56.355 43.333 ;
      RECT 53.831 43.231 56.401 43.287 ;
      RECT 53.877 43.185 56.447 43.241 ;
      RECT 53.923 43.139 56.493 43.195 ;
      RECT 53.969 43.093 56.539 43.149 ;
      RECT 54.015 43.047 56.585 43.103 ;
      RECT 54.061 43.001 56.631 43.057 ;
      RECT 54.107 42.955 56.677 43.011 ;
      RECT 54.153 42.909 56.723 42.965 ;
      RECT 54.199 42.863 56.769 42.919 ;
      RECT 54.245 42.817 56.815 42.873 ;
      RECT 54.291 42.771 56.861 42.827 ;
      RECT 54.337 42.725 56.907 42.781 ;
      RECT 54.383 42.679 56.953 42.735 ;
      RECT 54.429 42.633 56.999 42.689 ;
      RECT 54.475 42.587 57.045 42.643 ;
      RECT 54.521 42.541 57.091 42.597 ;
      RECT 54.567 42.495 57.137 42.551 ;
      RECT 54.613 42.449 57.183 42.505 ;
      RECT 54.659 42.403 57.229 42.459 ;
      RECT 54.705 42.357 57.275 42.413 ;
      RECT 54.751 42.311 57.321 42.367 ;
      RECT 54.797 42.265 57.367 42.321 ;
      RECT 54.843 42.219 57.413 42.275 ;
      RECT 54.889 42.173 57.459 42.229 ;
      RECT 54.935 42.127 57.505 42.183 ;
      RECT 54.981 42.081 57.551 42.137 ;
      RECT 55.027 42.035 57.597 42.091 ;
      RECT 55.073 41.989 57.643 42.045 ;
      RECT 55.119 41.943 57.689 41.999 ;
      RECT 55.165 41.897 57.735 41.953 ;
      RECT 55.211 41.851 57.781 41.907 ;
      RECT 55.257 41.805 57.827 41.861 ;
      RECT 55.303 41.759 57.873 41.815 ;
      RECT 55.349 41.713 57.919 41.769 ;
      RECT 55.395 41.667 57.965 41.723 ;
      RECT 55.441 41.621 58.011 41.677 ;
      RECT 55.487 41.575 58.057 41.631 ;
      RECT 55.533 41.529 58.103 41.585 ;
      RECT 55.579 41.483 58.149 41.539 ;
      RECT 55.625 41.437 58.195 41.493 ;
      RECT 55.671 41.391 58.241 41.447 ;
      RECT 55.717 41.345 58.287 41.401 ;
      RECT 55.763 41.299 58.333 41.355 ;
      RECT 55.809 41.253 58.379 41.309 ;
      RECT 55.855 41.207 58.425 41.263 ;
      RECT 55.901 41.161 58.471 41.217 ;
      RECT 55.947 41.115 58.517 41.171 ;
      RECT 55.993 41.069 58.563 41.125 ;
      RECT 56.039 41.023 58.609 41.079 ;
      RECT 56.085 40.977 58.655 41.033 ;
      RECT 56.131 40.931 58.701 40.987 ;
      RECT 56.177 40.885 58.747 40.941 ;
      RECT 56.223 40.839 58.793 40.895 ;
      RECT 56.269 40.793 58.839 40.849 ;
      RECT 56.315 40.747 58.885 40.803 ;
      RECT 56.361 40.701 58.931 40.757 ;
      RECT 56.407 40.655 58.977 40.711 ;
      RECT 56.453 40.609 59.023 40.665 ;
      RECT 56.499 40.563 59.069 40.619 ;
      RECT 56.545 40.517 59.115 40.573 ;
      RECT 56.591 40.471 59.161 40.527 ;
      RECT 56.637 40.425 59.207 40.481 ;
      RECT 56.683 40.379 59.253 40.435 ;
      RECT 56.729 40.333 59.299 40.389 ;
      RECT 56.775 40.287 59.345 40.343 ;
      RECT 56.821 40.241 59.391 40.297 ;
      RECT 56.867 40.195 59.437 40.251 ;
      RECT 56.913 40.149 59.483 40.205 ;
      RECT 56.959 40.103 59.529 40.159 ;
      RECT 57.005 40.057 59.575 40.113 ;
      RECT 57.051 40.011 59.621 40.067 ;
      RECT 57.097 39.965 59.667 40.021 ;
      RECT 57.143 39.919 59.713 39.975 ;
      RECT 57.189 39.873 59.759 39.929 ;
      RECT 57.235 39.827 59.805 39.883 ;
      RECT 57.281 39.781 59.851 39.837 ;
      RECT 57.327 39.735 59.897 39.791 ;
      RECT 57.373 39.689 59.943 39.745 ;
      RECT 57.419 39.643 59.989 39.699 ;
      RECT 57.465 39.597 60.035 39.653 ;
      RECT 57.511 39.551 60.081 39.607 ;
      RECT 57.557 39.505 60.127 39.561 ;
      RECT 57.603 39.459 60.173 39.515 ;
      RECT 57.649 39.413 60.219 39.469 ;
      RECT 57.695 39.367 60.265 39.423 ;
      RECT 57.741 39.321 60.311 39.377 ;
      RECT 57.787 39.275 60.357 39.331 ;
      RECT 57.833 39.229 60.403 39.285 ;
      RECT 57.879 39.183 60.449 39.239 ;
      RECT 57.925 39.137 60.495 39.193 ;
      RECT 57.971 39.091 60.541 39.147 ;
      RECT 58.017 39.045 60.587 39.101 ;
      RECT 58.063 38.999 60.633 39.055 ;
      RECT 58.109 38.953 60.679 39.009 ;
      RECT 58.155 38.907 60.725 38.963 ;
      RECT 58.201 38.861 60.771 38.917 ;
      RECT 58.247 38.815 60.817 38.871 ;
      RECT 58.293 38.769 60.863 38.825 ;
      RECT 58.339 38.723 60.909 38.779 ;
      RECT 58.385 38.677 60.955 38.733 ;
      RECT 58.431 38.631 61.001 38.687 ;
      RECT 58.477 38.585 61.047 38.641 ;
      RECT 58.523 38.539 61.093 38.595 ;
      RECT 58.569 38.493 61.139 38.549 ;
      RECT 58.615 38.447 61.185 38.503 ;
      RECT 58.661 38.401 61.231 38.457 ;
      RECT 58.707 38.355 61.277 38.411 ;
      RECT 58.753 38.309 61.323 38.365 ;
      RECT 58.799 38.263 61.369 38.319 ;
      RECT 58.845 38.217 61.415 38.273 ;
      RECT 58.891 38.171 61.461 38.227 ;
      RECT 58.937 38.125 61.507 38.181 ;
      RECT 58.983 38.079 61.553 38.135 ;
      RECT 59.029 38.033 61.599 38.089 ;
      RECT 59.075 37.987 61.645 38.043 ;
      RECT 59.121 37.941 61.691 37.997 ;
      RECT 59.167 37.895 61.737 37.951 ;
      RECT 59.213 37.849 61.783 37.905 ;
      RECT 59.259 37.803 61.829 37.859 ;
      RECT 59.305 37.757 61.875 37.813 ;
      RECT 59.351 37.711 61.921 37.767 ;
      RECT 59.397 37.665 61.967 37.721 ;
      RECT 59.443 37.619 62.013 37.675 ;
      RECT 59.489 37.573 62.059 37.629 ;
      RECT 59.535 37.527 62.105 37.583 ;
      RECT 59.581 37.481 62.151 37.537 ;
      RECT 59.627 37.435 62.197 37.491 ;
      RECT 59.673 37.389 62.243 37.445 ;
      RECT 59.719 37.343 62.289 37.399 ;
      RECT 59.765 37.297 62.335 37.353 ;
      RECT 59.811 37.251 62.381 37.307 ;
      RECT 59.857 37.205 62.427 37.261 ;
      RECT 59.903 37.159 62.473 37.215 ;
      RECT 59.949 37.113 62.519 37.169 ;
      RECT 59.995 37.067 62.565 37.123 ;
      RECT 60.041 37.021 62.611 37.077 ;
      RECT 60.087 36.975 62.657 37.031 ;
      RECT 60.133 36.929 62.703 36.985 ;
      RECT 60.179 36.883 62.749 36.939 ;
      RECT 60.225 36.837 62.795 36.893 ;
      RECT 60.271 36.791 62.841 36.847 ;
      RECT 60.317 36.745 62.887 36.801 ;
      RECT 60.363 36.699 62.933 36.755 ;
      RECT 60.409 36.653 62.979 36.709 ;
      RECT 62.939 34.146 62.979 36.709 ;
      RECT 60.455 36.607 63.025 36.663 ;
      RECT 62.94 34.122 63.025 36.663 ;
      RECT 60.501 36.561 63.071 36.617 ;
      RECT 62.986 34.076 63.071 36.617 ;
      RECT 60.547 36.515 63.117 36.571 ;
      RECT 63.032 34.03 63.117 36.571 ;
      RECT 60.593 36.469 63.163 36.525 ;
      RECT 63.078 33.984 63.163 36.525 ;
      RECT 60.639 36.423 63.209 36.479 ;
      RECT 63.124 33.938 63.209 36.479 ;
      RECT 60.685 36.377 63.255 36.433 ;
      RECT 63.17 33.892 63.255 36.433 ;
      RECT 60.731 36.331 63.301 36.387 ;
      RECT 63.216 33.846 63.301 36.387 ;
      RECT 60.777 36.285 63.347 36.341 ;
      RECT 63.262 33.8 63.347 36.341 ;
      RECT 60.823 36.239 63.393 36.295 ;
      RECT 63.308 33.754 63.393 36.295 ;
      RECT 60.869 36.193 63.439 36.249 ;
      RECT 63.354 33.708 63.439 36.249 ;
      RECT 60.915 36.147 63.485 36.203 ;
      RECT 63.4 33.662 63.485 36.203 ;
      RECT 60.961 36.101 63.531 36.157 ;
      RECT 63.446 33.616 63.531 36.157 ;
      RECT 61.007 36.055 63.577 36.111 ;
      RECT 63.492 33.57 63.577 36.111 ;
      RECT 61.053 36.009 63.623 36.065 ;
      RECT 63.538 33.524 63.623 36.065 ;
      RECT 61.099 35.963 63.669 36.019 ;
      RECT 63.584 33.478 63.669 36.019 ;
      RECT 61.145 35.917 63.715 35.973 ;
      RECT 63.63 33.432 63.715 35.973 ;
      RECT 61.191 35.871 63.761 35.927 ;
      RECT 63.676 33.386 63.761 35.927 ;
      RECT 61.237 35.825 63.807 35.881 ;
      RECT 63.722 33.34 63.807 35.881 ;
      RECT 61.283 35.779 63.853 35.835 ;
      RECT 63.768 33.294 63.853 35.835 ;
      RECT 61.329 35.733 63.899 35.789 ;
      RECT 63.814 33.248 63.899 35.789 ;
      RECT 61.375 35.687 63.945 35.743 ;
      RECT 63.86 33.202 63.945 35.743 ;
      RECT 61.421 35.641 63.991 35.697 ;
      RECT 63.906 33.156 63.991 35.697 ;
      RECT 61.467 35.595 64.037 35.651 ;
      RECT 63.952 33.11 64.037 35.651 ;
      RECT 61.513 35.549 64.083 35.605 ;
      RECT 63.998 33.064 64.083 35.605 ;
      RECT 61.559 35.503 64.129 35.559 ;
      RECT 64.044 33.018 64.129 35.559 ;
      RECT 61.605 35.457 64.175 35.513 ;
      RECT 64.09 32.972 64.175 35.513 ;
      RECT 61.651 35.411 64.221 35.467 ;
      RECT 64.136 32.926 64.221 35.467 ;
      RECT 61.697 35.365 64.267 35.421 ;
      RECT 64.182 32.88 64.267 35.421 ;
      RECT 61.743 35.319 64.313 35.375 ;
      RECT 64.228 32.834 64.313 35.375 ;
      RECT 61.789 35.273 64.359 35.329 ;
      RECT 64.274 32.788 64.359 35.329 ;
      RECT 61.835 35.227 64.405 35.283 ;
      RECT 64.32 32.742 64.405 35.283 ;
      RECT 61.881 35.181 64.451 35.237 ;
      RECT 64.366 32.696 64.451 35.237 ;
      RECT 61.927 35.135 64.497 35.191 ;
      RECT 64.412 32.65 64.497 35.191 ;
      RECT 61.973 35.089 64.543 35.145 ;
      RECT 64.458 32.604 64.543 35.145 ;
      RECT 62.019 35.043 64.589 35.099 ;
      RECT 64.504 32.558 64.589 35.099 ;
      RECT 62.065 34.997 64.635 35.053 ;
      RECT 64.55 32.512 64.635 35.053 ;
      RECT 62.111 34.951 64.681 35.007 ;
      RECT 64.596 32.466 64.681 35.007 ;
      RECT 62.157 34.905 64.727 34.961 ;
      RECT 64.642 32.42 64.727 34.961 ;
      RECT 62.203 34.859 64.773 34.915 ;
      RECT 64.688 32.374 64.773 34.915 ;
      RECT 62.249 34.813 64.819 34.869 ;
      RECT 64.734 32.328 64.819 34.869 ;
      RECT 62.295 34.767 64.865 34.823 ;
      RECT 64.78 32.282 64.865 34.823 ;
      RECT 62.341 34.721 64.911 34.777 ;
      RECT 64.826 32.236 64.911 34.777 ;
      RECT 62.387 34.675 64.957 34.731 ;
      RECT 64.872 32.19 64.957 34.731 ;
      RECT 62.433 34.629 65.003 34.685 ;
      RECT 64.918 32.144 65.003 34.685 ;
      RECT 62.479 34.583 65.049 34.639 ;
      RECT 64.964 32.098 65.049 34.639 ;
      RECT 62.525 34.537 65.095 34.593 ;
      RECT 65.01 32.052 65.095 34.593 ;
      RECT 62.571 34.491 65.141 34.547 ;
      RECT 65.056 32.006 65.141 34.547 ;
      RECT 62.617 34.445 65.187 34.501 ;
      RECT 65.102 31.96 65.187 34.501 ;
      RECT 62.663 34.399 65.233 34.455 ;
      RECT 65.148 31.914 65.233 34.455 ;
      RECT 62.709 34.353 65.279 34.409 ;
      RECT 65.194 31.868 65.279 34.409 ;
      RECT 62.755 34.307 65.325 34.363 ;
      RECT 65.24 31.822 65.325 34.363 ;
      RECT 62.801 34.261 65.371 34.317 ;
      RECT 65.286 31.776 65.371 34.317 ;
      RECT 62.847 34.215 65.417 34.271 ;
      RECT 65.332 31.73 65.417 34.271 ;
      RECT 62.893 34.169 65.463 34.225 ;
      RECT 65.378 31.684 65.463 34.225 ;
      RECT 65.424 31.638 65.509 34.179 ;
      RECT 65.47 31.592 65.555 34.133 ;
      RECT 65.516 31.546 65.601 34.087 ;
      RECT 65.562 31.5 65.647 34.041 ;
      RECT 65.608 31.454 65.693 33.995 ;
      RECT 65.654 31.408 65.739 33.949 ;
      RECT 65.7 31.362 65.785 33.903 ;
      RECT 65.746 31.316 65.831 33.857 ;
      RECT 65.792 31.27 65.877 33.811 ;
      RECT 65.838 31.224 65.923 33.765 ;
      RECT 65.884 31.178 65.969 33.719 ;
      RECT 65.93 31.132 66.015 33.673 ;
      RECT 65.976 31.086 66.061 33.627 ;
      RECT 66.022 31.04 66.107 33.581 ;
      RECT 66.068 30.994 66.153 33.535 ;
      RECT 66.114 30.948 66.199 33.489 ;
      RECT 66.16 30.902 66.245 33.443 ;
      RECT 66.206 30.856 66.291 33.397 ;
      RECT 66.252 30.81 66.337 33.351 ;
      RECT 66.298 30.764 66.383 33.305 ;
      RECT 66.344 30.718 66.429 33.259 ;
      RECT 66.39 30.672 66.475 33.213 ;
      RECT 66.436 30.626 66.521 33.167 ;
      RECT 66.482 30.58 66.567 33.121 ;
      RECT 66.528 30.534 66.613 33.075 ;
      RECT 66.574 30.488 66.659 33.029 ;
      RECT 66.62 30.442 66.705 32.983 ;
      RECT 66.666 30.396 66.751 32.937 ;
      RECT 66.712 30.35 66.797 32.891 ;
      RECT 66.758 30.304 66.843 32.845 ;
      RECT 66.804 30.258 66.889 32.799 ;
      RECT 66.85 30.212 66.935 32.753 ;
      RECT 66.896 30.166 66.981 32.707 ;
      RECT 66.942 30.12 67.027 32.661 ;
      RECT 66.988 30.074 67.073 32.615 ;
      RECT 67.034 30.028 67.119 32.569 ;
      RECT 67.08 29.982 67.165 32.523 ;
      RECT 67.126 29.936 67.211 32.477 ;
      RECT 67.172 29.89 67.257 32.431 ;
      RECT 67.218 29.844 67.303 32.385 ;
      RECT 67.264 29.798 67.349 32.339 ;
      RECT 67.31 29.752 67.395 32.293 ;
      RECT 67.356 29.706 67.441 32.247 ;
      RECT 67.402 29.66 67.487 32.201 ;
      RECT 67.448 29.614 67.533 32.155 ;
      RECT 67.494 29.568 67.579 32.109 ;
      RECT 67.54 29.522 67.625 32.063 ;
      RECT 67.586 29.476 67.671 32.017 ;
      RECT 67.632 29.43 67.717 31.971 ;
      RECT 67.678 29.384 67.763 31.925 ;
      RECT 67.724 29.338 67.809 31.879 ;
      RECT 67.77 29.292 67.855 31.833 ;
      RECT 67.816 29.246 67.901 31.787 ;
      RECT 67.862 29.199 67.947 31.741 ;
      RECT 67.908 29.175 67.993 31.695 ;
      RECT 67.908 29.175 68.039 31.649 ;
      RECT 67.908 29.175 68.085 31.603 ;
      RECT 67.908 29.175 68.131 31.557 ;
      RECT 67.908 29.175 68.177 31.511 ;
      RECT 67.908 29.175 68.223 31.465 ;
      RECT 67.908 29.175 68.269 31.419 ;
      RECT 67.908 29.175 68.315 31.373 ;
      RECT 67.908 29.175 68.361 31.327 ;
      RECT 67.908 29.175 68.407 31.281 ;
      RECT 67.908 29.175 68.453 31.235 ;
      RECT 67.908 29.175 68.499 31.189 ;
      RECT 67.908 29.175 68.545 31.143 ;
      RECT 67.908 29.175 68.591 31.097 ;
      RECT 67.908 29.175 68.637 31.051 ;
      RECT 67.908 29.175 68.683 31.005 ;
      RECT 67.908 29.175 68.729 30.959 ;
      RECT 67.908 29.175 68.775 30.913 ;
      RECT 67.908 29.175 68.821 30.867 ;
      RECT 67.908 29.175 68.867 30.821 ;
      RECT 67.908 29.175 68.913 30.775 ;
      RECT 67.908 29.175 68.959 30.729 ;
      RECT 67.908 29.175 69.005 30.683 ;
      RECT 67.908 29.175 69.051 30.637 ;
      RECT 67.908 29.175 69.097 30.591 ;
      RECT 67.908 29.175 69.143 30.545 ;
      RECT 67.908 29.175 69.189 30.499 ;
      RECT 67.908 29.175 69.235 30.453 ;
      RECT 67.908 29.175 69.281 30.407 ;
      RECT 67.908 29.175 69.327 30.361 ;
      RECT 66.758 30.304 69.34 30.331 ;
      RECT 67.908 29.175 110 30.325 ;
      RECT 42.675 74.637 43.825 110 ;
      RECT 42.675 74.637 43.871 76.067 ;
      RECT 42.675 74.637 43.917 76.021 ;
      RECT 42.675 74.637 43.963 75.975 ;
      RECT 42.675 74.637 44.009 75.929 ;
      RECT 42.675 74.637 44.055 75.883 ;
      RECT 42.675 74.637 44.101 75.837 ;
      RECT 42.675 74.637 44.147 75.791 ;
      RECT 42.675 74.637 44.193 75.745 ;
      RECT 42.675 74.637 44.239 75.699 ;
      RECT 42.675 74.637 44.285 75.653 ;
      RECT 42.675 74.637 44.331 75.607 ;
      RECT 42.675 74.637 44.377 75.561 ;
      RECT 42.675 74.637 44.423 75.515 ;
      RECT 42.675 74.637 44.469 75.469 ;
      RECT 42.675 74.637 44.515 75.423 ;
      RECT 42.675 74.637 44.561 75.377 ;
      RECT 42.675 74.637 44.607 75.331 ;
      RECT 42.675 74.637 44.653 75.285 ;
      RECT 42.675 74.637 44.699 75.239 ;
      RECT 42.675 74.637 44.745 75.193 ;
      RECT 42.675 74.637 44.791 75.147 ;
      RECT 42.675 74.637 44.837 75.101 ;
      RECT 42.675 74.637 44.883 75.055 ;
      RECT 42.675 74.637 44.929 75.009 ;
      RECT 42.675 74.637 44.975 74.963 ;
      RECT 42.675 74.637 45.021 74.917 ;
      RECT 42.675 74.637 45.067 74.871 ;
      RECT 42.675 74.637 45.113 74.825 ;
      RECT 42.675 74.637 45.159 74.779 ;
      RECT 42.675 74.637 45.205 74.733 ;
      RECT 42.675 74.637 45.251 74.687 ;
      RECT 42.721 74.591 45.297 74.641 ;
      RECT 42.767 74.545 45.343 74.595 ;
      RECT 42.813 74.499 45.389 74.549 ;
      RECT 42.859 74.453 45.435 74.503 ;
      RECT 42.905 74.407 45.481 74.457 ;
      RECT 42.951 74.361 45.527 74.411 ;
      RECT 42.997 74.315 45.573 74.365 ;
      RECT 43.043 74.269 45.619 74.319 ;
      RECT 43.089 74.223 45.665 74.273 ;
      RECT 43.135 74.177 45.711 74.227 ;
      RECT 43.181 74.131 45.757 74.181 ;
      RECT 43.227 74.085 45.803 74.135 ;
      RECT 43.273 74.039 45.849 74.089 ;
      RECT 43.319 73.993 45.895 74.043 ;
      RECT 43.365 73.947 45.941 73.997 ;
      RECT 43.411 73.901 45.987 73.951 ;
      RECT 43.457 73.855 46.033 73.905 ;
      RECT 43.503 73.809 46.079 73.859 ;
      RECT 43.549 73.763 46.125 73.813 ;
      RECT 43.595 73.717 46.171 73.767 ;
      RECT 43.641 73.671 46.217 73.721 ;
      RECT 43.687 73.625 46.263 73.675 ;
      RECT 43.733 73.579 46.309 73.629 ;
      RECT 43.779 73.533 46.355 73.583 ;
      RECT 43.825 73.487 46.401 73.537 ;
      RECT 43.871 73.441 46.447 73.491 ;
      RECT 43.917 73.395 46.493 73.445 ;
      RECT 43.963 73.349 46.539 73.399 ;
      RECT 44.009 73.303 46.585 73.353 ;
      RECT 44.055 73.257 46.631 73.307 ;
      RECT 44.101 73.211 46.677 73.261 ;
      RECT 44.147 73.165 46.723 73.215 ;
      RECT 44.193 73.119 46.769 73.169 ;
      RECT 44.239 73.073 46.815 73.123 ;
      RECT 44.285 73.027 46.861 73.077 ;
      RECT 44.331 72.981 46.907 73.031 ;
      RECT 44.377 72.935 46.953 72.985 ;
      RECT 44.423 72.889 46.999 72.939 ;
      RECT 44.469 72.843 47.045 72.893 ;
      RECT 44.515 72.797 47.091 72.847 ;
      RECT 44.561 72.751 47.137 72.801 ;
      RECT 44.607 72.705 47.183 72.755 ;
      RECT 44.653 72.659 47.229 72.709 ;
      RECT 44.699 72.613 47.275 72.663 ;
      RECT 44.745 72.567 47.321 72.617 ;
      RECT 44.791 72.521 47.367 72.571 ;
      RECT 44.837 72.475 47.413 72.525 ;
      RECT 44.883 72.429 47.459 72.479 ;
      RECT 44.929 72.383 47.505 72.433 ;
      RECT 44.975 72.337 47.551 72.387 ;
      RECT 45.021 72.291 47.597 72.341 ;
      RECT 45.067 72.245 47.643 72.295 ;
      RECT 45.113 72.199 47.689 72.249 ;
      RECT 45.159 72.153 47.735 72.203 ;
      RECT 45.205 72.107 47.781 72.157 ;
      RECT 45.251 72.061 47.827 72.111 ;
      RECT 45.297 72.015 47.873 72.065 ;
      RECT 45.343 71.969 47.919 72.019 ;
      RECT 45.389 71.923 47.965 71.973 ;
      RECT 45.435 71.877 48.011 71.927 ;
      RECT 45.481 71.831 48.057 71.881 ;
      RECT 45.527 71.785 48.103 71.835 ;
      RECT 45.573 71.739 48.149 71.789 ;
      RECT 45.619 71.693 48.195 71.743 ;
      RECT 45.665 71.647 48.241 71.697 ;
      RECT 45.711 71.601 48.287 71.651 ;
      RECT 45.757 71.555 48.333 71.605 ;
      RECT 45.803 71.509 48.379 71.559 ;
      RECT 45.849 71.463 48.425 71.513 ;
      RECT 45.895 71.417 48.471 71.467 ;
      RECT 45.941 71.371 48.517 71.421 ;
      RECT 45.987 71.325 48.563 71.375 ;
      RECT 46.033 71.279 48.609 71.329 ;
      RECT 46.079 71.233 48.655 71.283 ;
      RECT 46.125 71.187 48.701 71.237 ;
      RECT 46.171 71.141 48.747 71.191 ;
      RECT 46.217 71.095 48.793 71.145 ;
      RECT 46.263 71.049 48.839 71.099 ;
      RECT 46.309 71.003 48.885 71.053 ;
      RECT 46.355 70.957 48.931 71.007 ;
      RECT 46.401 70.911 48.977 70.961 ;
      RECT 46.447 70.865 49.023 70.915 ;
      RECT 46.493 70.819 49.069 70.869 ;
      RECT 46.539 70.773 49.115 70.823 ;
      RECT 46.585 70.727 49.161 70.777 ;
      RECT 46.631 70.681 49.207 70.731 ;
      RECT 46.677 70.635 49.253 70.685 ;
      RECT 46.723 70.589 49.299 70.639 ;
      RECT 46.769 70.543 49.345 70.593 ;
      RECT 46.815 70.497 49.391 70.547 ;
      RECT 46.861 70.451 49.437 70.501 ;
      RECT 46.907 70.405 49.483 70.455 ;
      RECT 46.953 70.359 49.529 70.409 ;
      RECT 46.999 70.313 49.575 70.363 ;
      RECT 47.045 70.267 49.621 70.317 ;
      RECT 47.091 70.221 49.667 70.271 ;
      RECT 47.137 70.175 49.713 70.225 ;
      RECT 47.183 70.129 49.759 70.179 ;
      RECT 47.229 70.083 49.805 70.133 ;
      RECT 47.275 70.037 49.851 70.087 ;
      RECT 47.321 69.991 49.897 70.041 ;
      RECT 47.367 69.945 49.943 69.995 ;
      RECT 47.413 69.899 49.989 69.949 ;
      RECT 47.459 69.853 50.035 69.903 ;
      RECT 47.505 69.807 50.081 69.857 ;
      RECT 47.551 69.761 50.127 69.811 ;
      RECT 47.597 69.715 50.173 69.765 ;
      RECT 47.643 69.669 50.219 69.719 ;
      RECT 47.689 69.623 50.265 69.673 ;
      RECT 47.735 69.577 50.311 69.627 ;
      RECT 47.781 69.531 50.357 69.581 ;
      RECT 47.827 69.485 50.403 69.535 ;
      RECT 47.873 69.439 50.449 69.489 ;
      RECT 47.919 69.393 50.495 69.443 ;
      RECT 47.965 69.347 50.541 69.397 ;
      RECT 48.011 69.301 50.587 69.351 ;
      RECT 48.057 69.255 50.633 69.305 ;
      RECT 48.103 69.209 50.679 69.259 ;
      RECT 48.149 69.163 50.725 69.213 ;
      RECT 48.195 69.117 50.771 69.167 ;
      RECT 48.241 69.071 50.817 69.121 ;
      RECT 48.287 69.025 50.863 69.075 ;
      RECT 48.333 68.979 50.909 69.029 ;
      RECT 48.379 68.933 50.955 68.983 ;
      RECT 48.425 68.887 51.001 68.937 ;
      RECT 48.471 68.841 51.047 68.891 ;
      RECT 48.517 68.795 51.093 68.845 ;
      RECT 48.563 68.749 51.139 68.799 ;
      RECT 48.609 68.703 51.185 68.753 ;
      RECT 48.655 68.657 51.231 68.707 ;
      RECT 48.701 68.611 51.277 68.661 ;
      RECT 48.747 68.565 51.323 68.615 ;
      RECT 48.793 68.519 51.369 68.569 ;
      RECT 48.839 68.473 51.415 68.523 ;
      RECT 48.885 68.427 51.461 68.477 ;
      RECT 48.931 68.381 51.507 68.431 ;
      RECT 48.977 68.335 51.553 68.385 ;
      RECT 49.023 68.289 51.599 68.339 ;
      RECT 49.069 68.243 51.645 68.293 ;
      RECT 49.115 68.197 51.691 68.247 ;
      RECT 49.161 68.151 51.737 68.201 ;
      RECT 49.207 68.105 51.783 68.155 ;
      RECT 49.253 68.059 51.829 68.109 ;
      RECT 49.299 68.013 51.875 68.063 ;
      RECT 49.345 67.967 51.921 68.017 ;
      RECT 49.391 67.921 51.967 67.971 ;
      RECT 49.437 67.875 52.013 67.925 ;
      RECT 49.483 67.829 52.059 67.879 ;
      RECT 49.529 67.783 52.105 67.833 ;
      RECT 49.575 67.737 52.151 67.787 ;
      RECT 49.621 67.691 52.197 67.741 ;
      RECT 49.667 67.645 52.243 67.695 ;
      RECT 49.713 67.599 52.289 67.649 ;
      RECT 49.759 67.553 52.335 67.603 ;
      RECT 49.805 67.507 52.381 67.557 ;
      RECT 49.851 67.461 52.427 67.511 ;
      RECT 49.897 67.415 52.473 67.465 ;
      RECT 49.943 67.369 52.519 67.419 ;
      RECT 49.989 67.323 52.565 67.373 ;
      RECT 50.035 67.277 52.611 67.327 ;
      RECT 50.081 67.231 52.657 67.281 ;
      RECT 50.127 67.185 52.703 67.235 ;
      RECT 50.173 67.139 52.749 67.189 ;
      RECT 50.219 67.093 52.795 67.143 ;
      RECT 50.265 67.047 52.841 67.097 ;
      RECT 50.311 67.001 52.887 67.051 ;
      RECT 50.357 66.955 52.933 67.005 ;
      RECT 50.403 66.909 52.979 66.959 ;
      RECT 50.449 66.863 53.025 66.913 ;
      RECT 50.495 66.817 53.071 66.867 ;
      RECT 50.541 66.771 53.117 66.821 ;
      RECT 50.587 66.725 53.163 66.775 ;
      RECT 50.633 66.679 53.209 66.729 ;
      RECT 50.679 66.633 53.255 66.683 ;
      RECT 50.725 66.587 53.301 66.637 ;
      RECT 50.771 66.541 53.347 66.591 ;
      RECT 50.817 66.495 53.393 66.545 ;
      RECT 50.863 66.449 53.439 66.499 ;
      RECT 50.909 66.403 53.485 66.453 ;
      RECT 50.955 66.357 53.531 66.407 ;
      RECT 51.001 66.311 53.577 66.361 ;
      RECT 51.047 66.265 53.623 66.315 ;
      RECT 51.093 66.219 53.669 66.269 ;
      RECT 51.139 66.173 53.715 66.223 ;
      RECT 51.185 66.127 53.761 66.177 ;
      RECT 51.231 66.081 53.807 66.131 ;
      RECT 51.277 66.035 53.853 66.085 ;
      RECT 51.323 65.989 53.899 66.039 ;
      RECT 51.369 65.943 53.945 65.993 ;
      RECT 51.415 65.897 53.991 65.947 ;
      RECT 51.461 65.851 54.037 65.901 ;
      RECT 51.507 65.805 54.083 65.855 ;
      RECT 51.553 65.759 54.129 65.809 ;
      RECT 51.599 65.713 54.175 65.763 ;
      RECT 51.645 65.667 54.221 65.717 ;
      RECT 51.691 65.621 54.267 65.671 ;
      RECT 51.737 65.575 54.313 65.625 ;
      RECT 51.783 65.529 54.359 65.579 ;
      RECT 51.829 65.483 54.405 65.533 ;
      RECT 51.875 65.437 54.451 65.487 ;
      RECT 51.921 65.391 54.497 65.441 ;
      RECT 51.967 65.345 54.543 65.395 ;
      RECT 52.013 65.299 54.589 65.349 ;
      RECT 52.059 65.253 54.635 65.303 ;
      RECT 52.105 65.207 54.681 65.257 ;
      RECT 52.151 65.161 54.727 65.211 ;
      RECT 52.197 65.115 54.773 65.165 ;
      RECT 52.243 65.069 54.819 65.119 ;
      RECT 52.289 65.023 54.865 65.073 ;
      RECT 52.335 64.977 54.911 65.027 ;
      RECT 52.381 64.931 54.957 64.981 ;
      RECT 52.427 64.885 55.003 64.935 ;
      RECT 52.473 64.839 55.049 64.889 ;
      RECT 52.519 64.793 55.095 64.843 ;
      RECT 52.565 64.747 55.141 64.797 ;
      RECT 52.611 64.701 55.187 64.751 ;
      RECT 52.657 64.655 55.233 64.705 ;
      RECT 52.703 64.609 55.279 64.659 ;
      RECT 52.749 64.563 55.325 64.613 ;
      RECT 52.795 64.517 55.371 64.567 ;
      RECT 52.841 64.471 55.417 64.521 ;
      RECT 52.887 64.425 55.463 64.475 ;
      RECT 52.933 64.379 55.509 64.429 ;
      RECT 52.979 64.333 55.555 64.383 ;
      RECT 53.025 64.287 55.601 64.337 ;
      RECT 53.071 64.241 55.647 64.291 ;
      RECT 53.117 64.195 55.693 64.245 ;
      RECT 53.163 64.149 55.739 64.199 ;
      RECT 53.209 64.103 55.785 64.153 ;
      RECT 53.255 64.057 55.825 64.11 ;
      RECT 53.301 64.011 55.871 64.067 ;
      RECT 53.347 63.965 55.917 64.021 ;
      RECT 53.393 63.919 55.963 63.975 ;
      RECT 53.439 63.873 56.009 63.929 ;
      RECT 53.485 63.827 56.055 63.883 ;
      RECT 53.531 63.781 56.101 63.837 ;
      RECT 53.577 63.735 56.147 63.791 ;
      RECT 53.623 63.689 56.193 63.745 ;
      RECT 53.669 63.643 56.239 63.699 ;
      RECT 53.715 63.597 56.285 63.653 ;
      RECT 53.761 63.551 56.331 63.607 ;
      RECT 53.807 63.505 56.377 63.561 ;
      RECT 53.853 63.459 56.423 63.515 ;
      RECT 53.899 63.413 56.469 63.469 ;
      RECT 53.945 63.367 56.515 63.423 ;
      RECT 53.991 63.321 56.561 63.377 ;
      RECT 54.037 63.275 56.607 63.331 ;
      RECT 54.083 63.229 56.653 63.285 ;
      RECT 54.129 63.183 56.699 63.239 ;
      RECT 54.175 63.137 56.745 63.193 ;
      RECT 54.221 63.091 56.791 63.147 ;
      RECT 54.267 63.045 56.837 63.101 ;
      RECT 54.313 62.999 56.883 63.055 ;
      RECT 54.359 62.953 56.929 63.009 ;
      RECT 54.405 62.907 56.975 62.963 ;
      RECT 54.451 62.861 57.021 62.917 ;
      RECT 54.497 62.815 57.067 62.871 ;
      RECT 54.543 62.769 57.113 62.825 ;
      RECT 54.589 62.723 57.159 62.779 ;
      RECT 54.635 62.677 57.205 62.733 ;
      RECT 54.681 62.631 57.251 62.687 ;
      RECT 54.727 62.585 57.297 62.641 ;
      RECT 54.773 62.539 57.343 62.595 ;
      RECT 54.819 62.493 57.389 62.549 ;
      RECT 54.865 62.447 57.435 62.503 ;
      RECT 54.911 62.401 57.481 62.457 ;
      RECT 54.957 62.355 57.527 62.411 ;
      RECT 55.003 62.309 57.573 62.365 ;
      RECT 55.049 62.263 57.619 62.319 ;
      RECT 55.095 62.217 57.665 62.273 ;
      RECT 55.141 62.171 57.711 62.227 ;
      RECT 55.187 62.125 57.757 62.181 ;
      RECT 55.233 62.079 57.803 62.135 ;
      RECT 55.279 62.033 57.849 62.089 ;
      RECT 55.325 61.987 57.895 62.043 ;
      RECT 55.371 61.941 57.941 61.997 ;
      RECT 55.417 61.895 57.987 61.951 ;
      RECT 55.463 61.849 58.033 61.905 ;
      RECT 55.509 61.803 58.079 61.859 ;
      RECT 55.555 61.757 58.125 61.813 ;
      RECT 55.601 61.711 58.171 61.767 ;
      RECT 55.647 61.665 58.217 61.721 ;
      RECT 55.693 61.619 58.263 61.675 ;
      RECT 55.739 61.573 58.309 61.629 ;
      RECT 55.785 61.527 58.355 61.583 ;
      RECT 55.831 61.481 58.401 61.537 ;
      RECT 55.877 61.435 58.447 61.491 ;
      RECT 55.923 61.389 58.493 61.445 ;
      RECT 55.969 61.343 58.539 61.399 ;
      RECT 56.015 61.297 58.585 61.353 ;
      RECT 56.061 61.251 58.631 61.307 ;
      RECT 56.107 61.205 58.677 61.261 ;
      RECT 56.153 61.159 58.723 61.215 ;
      RECT 56.199 61.113 58.769 61.169 ;
      RECT 56.245 61.067 58.815 61.123 ;
      RECT 56.291 61.021 58.861 61.077 ;
      RECT 56.337 60.975 58.907 61.031 ;
      RECT 56.383 60.929 58.953 60.985 ;
      RECT 56.429 60.883 58.999 60.939 ;
      RECT 56.475 60.837 59.045 60.893 ;
      RECT 56.521 60.791 59.091 60.847 ;
      RECT 56.567 60.745 59.137 60.801 ;
      RECT 56.613 60.699 59.183 60.755 ;
      RECT 56.659 60.653 59.229 60.709 ;
      RECT 56.705 60.607 59.275 60.663 ;
      RECT 56.751 60.561 59.321 60.617 ;
      RECT 56.797 60.515 59.367 60.571 ;
      RECT 56.843 60.469 59.413 60.525 ;
      RECT 56.889 60.423 59.459 60.479 ;
      RECT 56.935 60.377 59.505 60.433 ;
      RECT 56.981 60.331 59.551 60.387 ;
      RECT 57.027 60.285 59.597 60.341 ;
      RECT 57.073 60.239 59.643 60.295 ;
      RECT 57.119 60.193 59.689 60.249 ;
      RECT 57.165 60.147 59.735 60.203 ;
      RECT 57.211 60.101 59.781 60.157 ;
      RECT 57.257 60.055 59.827 60.111 ;
      RECT 57.303 60.009 59.873 60.065 ;
      RECT 57.349 59.963 59.919 60.019 ;
      RECT 57.395 59.917 59.965 59.973 ;
      RECT 57.441 59.871 60.011 59.927 ;
      RECT 57.487 59.825 60.057 59.881 ;
      RECT 57.533 59.779 60.103 59.835 ;
      RECT 57.579 59.733 60.149 59.789 ;
      RECT 57.625 59.687 60.195 59.743 ;
      RECT 57.671 59.641 60.241 59.697 ;
      RECT 57.717 59.595 60.287 59.651 ;
      RECT 57.763 59.549 60.333 59.605 ;
      RECT 57.809 59.503 60.379 59.559 ;
      RECT 57.855 59.457 60.425 59.513 ;
      RECT 57.901 59.411 60.471 59.467 ;
      RECT 57.947 59.365 60.517 59.421 ;
      RECT 57.993 59.319 60.563 59.375 ;
      RECT 58.039 59.273 60.609 59.329 ;
      RECT 58.085 59.227 60.655 59.283 ;
      RECT 58.131 59.181 60.701 59.237 ;
      RECT 58.177 59.135 60.747 59.191 ;
      RECT 58.223 59.089 60.793 59.145 ;
      RECT 58.269 59.043 60.839 59.099 ;
      RECT 58.315 58.997 60.885 59.053 ;
      RECT 58.361 58.951 60.931 59.007 ;
      RECT 58.407 58.905 60.977 58.961 ;
      RECT 58.453 58.859 61.023 58.915 ;
      RECT 58.499 58.813 61.069 58.869 ;
      RECT 58.545 58.767 61.115 58.823 ;
      RECT 58.591 58.721 61.161 58.777 ;
      RECT 58.637 58.675 61.207 58.731 ;
      RECT 58.683 58.629 61.253 58.685 ;
      RECT 58.729 58.583 61.299 58.639 ;
      RECT 58.775 58.537 61.345 58.593 ;
      RECT 58.821 58.491 61.391 58.547 ;
      RECT 58.867 58.445 61.437 58.501 ;
      RECT 58.913 58.399 61.483 58.455 ;
      RECT 58.959 58.353 61.529 58.409 ;
      RECT 59.005 58.307 61.575 58.363 ;
      RECT 59.051 58.261 61.621 58.317 ;
      RECT 59.097 58.215 61.667 58.271 ;
      RECT 59.143 58.169 61.713 58.225 ;
      RECT 59.189 58.123 61.759 58.179 ;
      RECT 59.235 58.077 61.805 58.133 ;
      RECT 59.281 58.031 61.851 58.087 ;
      RECT 59.327 57.985 61.897 58.041 ;
      RECT 59.373 57.939 61.943 57.995 ;
      RECT 59.419 57.893 61.989 57.949 ;
      RECT 59.465 57.847 62.035 57.903 ;
      RECT 59.511 57.801 62.081 57.857 ;
      RECT 59.557 57.755 62.127 57.811 ;
      RECT 59.603 57.709 62.173 57.765 ;
      RECT 59.649 57.663 62.219 57.719 ;
      RECT 59.695 57.617 62.265 57.673 ;
      RECT 59.741 57.571 62.311 57.627 ;
      RECT 59.787 57.525 62.357 57.581 ;
      RECT 59.833 57.479 62.403 57.535 ;
      RECT 59.879 57.433 62.449 57.489 ;
      RECT 59.925 57.387 62.495 57.443 ;
      RECT 59.971 57.341 62.541 57.397 ;
      RECT 60.017 57.295 62.587 57.351 ;
      RECT 60.063 57.249 62.633 57.305 ;
      RECT 60.109 57.203 62.679 57.259 ;
      RECT 60.155 57.157 62.725 57.213 ;
      RECT 60.201 57.111 62.771 57.167 ;
      RECT 60.247 57.065 62.817 57.121 ;
      RECT 60.293 57.019 62.863 57.075 ;
      RECT 60.339 56.973 62.909 57.029 ;
      RECT 60.385 56.927 62.955 56.983 ;
      RECT 60.431 56.881 63.001 56.937 ;
      RECT 60.477 56.835 63.047 56.891 ;
      RECT 60.523 56.789 63.093 56.845 ;
      RECT 60.569 56.743 63.139 56.799 ;
      RECT 60.615 56.697 63.185 56.753 ;
      RECT 60.661 56.651 63.231 56.707 ;
      RECT 60.707 56.605 63.277 56.661 ;
      RECT 60.753 56.559 63.323 56.615 ;
      RECT 60.799 56.513 63.369 56.569 ;
      RECT 60.845 56.467 63.415 56.523 ;
      RECT 60.891 56.421 63.461 56.477 ;
      RECT 60.937 56.375 63.507 56.431 ;
      RECT 60.983 56.329 63.553 56.385 ;
      RECT 61.029 56.283 63.599 56.339 ;
      RECT 61.075 56.237 63.645 56.293 ;
      RECT 61.121 56.191 63.691 56.247 ;
      RECT 61.167 56.145 63.737 56.201 ;
      RECT 61.213 56.099 63.783 56.155 ;
      RECT 61.259 56.053 63.829 56.109 ;
      RECT 61.305 56.007 63.875 56.063 ;
      RECT 61.351 55.961 63.921 56.017 ;
      RECT 61.397 55.915 63.967 55.971 ;
      RECT 61.443 55.869 64.013 55.925 ;
      RECT 61.489 55.823 64.059 55.879 ;
      RECT 61.535 55.777 64.105 55.833 ;
      RECT 61.581 55.731 64.151 55.787 ;
      RECT 61.627 55.685 64.197 55.741 ;
      RECT 61.673 55.639 64.243 55.695 ;
      RECT 61.719 55.593 64.289 55.649 ;
      RECT 61.765 55.547 64.335 55.603 ;
      RECT 61.811 55.501 64.381 55.557 ;
      RECT 61.857 55.455 64.427 55.511 ;
      RECT 61.903 55.409 64.473 55.465 ;
      RECT 61.949 55.363 64.519 55.419 ;
      RECT 61.995 55.317 64.565 55.373 ;
      RECT 62.041 55.271 64.611 55.327 ;
      RECT 62.087 55.225 64.657 55.281 ;
      RECT 62.133 55.179 64.703 55.235 ;
      RECT 62.179 55.133 64.749 55.189 ;
      RECT 62.225 55.087 64.795 55.143 ;
      RECT 62.271 55.041 64.841 55.097 ;
      RECT 62.317 54.995 64.887 55.051 ;
      RECT 62.363 54.949 64.933 55.005 ;
      RECT 62.409 54.903 64.979 54.959 ;
      RECT 62.455 54.857 65.025 54.913 ;
      RECT 62.501 54.811 65.071 54.867 ;
      RECT 62.547 54.765 65.117 54.821 ;
      RECT 62.593 54.719 65.163 54.775 ;
      RECT 62.639 54.673 65.209 54.729 ;
      RECT 62.685 54.627 65.255 54.683 ;
      RECT 62.731 54.581 65.301 54.637 ;
      RECT 62.777 54.535 65.347 54.591 ;
      RECT 62.823 54.489 65.393 54.545 ;
      RECT 62.869 54.443 65.439 54.499 ;
      RECT 62.915 54.397 65.485 54.453 ;
      RECT 62.961 54.351 65.531 54.407 ;
      RECT 63.007 54.305 65.577 54.361 ;
      RECT 63.053 54.259 65.623 54.315 ;
      RECT 63.099 54.213 65.669 54.269 ;
      RECT 63.145 54.167 65.715 54.223 ;
      RECT 63.191 54.121 65.761 54.177 ;
      RECT 63.237 54.075 65.807 54.131 ;
      RECT 63.283 54.029 65.853 54.085 ;
      RECT 63.329 53.983 65.899 54.039 ;
      RECT 63.375 53.937 65.945 53.993 ;
      RECT 63.421 53.891 65.991 53.947 ;
      RECT 63.467 53.845 66.037 53.901 ;
      RECT 63.513 53.799 66.083 53.855 ;
      RECT 63.559 53.753 66.129 53.809 ;
      RECT 63.605 53.707 66.175 53.763 ;
      RECT 63.651 53.661 66.221 53.717 ;
      RECT 63.697 53.615 66.267 53.671 ;
      RECT 63.743 53.569 66.313 53.625 ;
      RECT 63.789 53.523 66.359 53.579 ;
      RECT 63.835 53.477 66.405 53.533 ;
      RECT 63.881 53.431 66.451 53.487 ;
      RECT 63.927 53.385 66.497 53.441 ;
      RECT 63.973 53.339 66.543 53.395 ;
      RECT 64.019 53.293 66.589 53.349 ;
      RECT 64.065 53.247 66.635 53.303 ;
      RECT 64.111 53.201 66.681 53.257 ;
      RECT 64.157 53.155 66.727 53.211 ;
      RECT 64.203 53.109 66.773 53.165 ;
      RECT 64.249 53.063 66.819 53.119 ;
      RECT 64.295 53.017 66.865 53.073 ;
      RECT 64.341 52.971 66.911 53.027 ;
      RECT 64.387 52.925 66.957 52.981 ;
      RECT 64.433 52.879 67.003 52.935 ;
      RECT 64.479 52.833 67.049 52.889 ;
      RECT 64.525 52.787 67.095 52.843 ;
      RECT 64.571 52.741 67.141 52.797 ;
      RECT 64.617 52.695 67.187 52.751 ;
      RECT 64.663 52.649 67.233 52.705 ;
      RECT 64.709 52.603 67.279 52.659 ;
      RECT 64.755 52.557 67.325 52.613 ;
      RECT 64.801 52.511 67.371 52.567 ;
      RECT 64.847 52.465 67.417 52.521 ;
      RECT 64.893 52.419 67.463 52.475 ;
      RECT 64.939 52.373 67.509 52.429 ;
      RECT 64.985 52.327 67.555 52.383 ;
      RECT 65.031 52.281 67.601 52.337 ;
      RECT 65.077 52.235 67.647 52.291 ;
      RECT 65.123 52.189 67.693 52.245 ;
      RECT 65.169 52.143 67.739 52.199 ;
      RECT 65.215 52.097 67.785 52.153 ;
      RECT 65.261 52.051 67.831 52.107 ;
      RECT 65.307 52.005 67.877 52.061 ;
      RECT 65.353 51.959 67.923 52.015 ;
      RECT 65.399 51.913 67.969 51.969 ;
      RECT 65.445 51.867 68.015 51.923 ;
      RECT 65.491 51.821 68.061 51.877 ;
      RECT 65.537 51.775 68.107 51.831 ;
      RECT 65.583 51.729 68.153 51.785 ;
      RECT 65.629 51.683 68.199 51.739 ;
      RECT 65.675 51.637 68.245 51.693 ;
      RECT 65.721 51.591 68.291 51.647 ;
      RECT 65.767 51.545 68.337 51.601 ;
      RECT 65.813 51.499 68.383 51.555 ;
      RECT 65.859 51.453 68.429 51.509 ;
      RECT 65.905 51.407 68.475 51.463 ;
      RECT 65.951 51.361 68.521 51.417 ;
      RECT 65.997 51.315 68.567 51.371 ;
      RECT 66.043 51.269 68.613 51.325 ;
      RECT 66.089 51.223 68.659 51.279 ;
      RECT 66.135 51.177 68.705 51.233 ;
      RECT 66.181 51.131 68.751 51.187 ;
      RECT 66.227 51.085 68.797 51.141 ;
      RECT 66.273 51.039 68.843 51.095 ;
      RECT 66.319 50.993 68.889 51.049 ;
      RECT 66.365 50.947 68.935 51.003 ;
      RECT 66.411 50.901 68.981 50.957 ;
      RECT 66.457 50.855 69.027 50.911 ;
      RECT 66.503 50.809 69.073 50.865 ;
      RECT 66.549 50.763 69.119 50.819 ;
      RECT 66.595 50.717 69.165 50.773 ;
      RECT 66.641 50.671 69.211 50.727 ;
      RECT 66.687 50.625 69.257 50.681 ;
      RECT 66.733 50.579 69.303 50.635 ;
      RECT 66.779 50.533 69.349 50.589 ;
      RECT 66.825 50.487 69.395 50.543 ;
      RECT 66.871 50.441 69.441 50.497 ;
      RECT 66.917 50.395 69.487 50.451 ;
      RECT 66.963 50.349 69.533 50.405 ;
      RECT 67.009 50.303 69.579 50.359 ;
      RECT 67.055 50.257 69.625 50.313 ;
      RECT 67.101 50.211 69.671 50.267 ;
      RECT 67.147 50.165 69.717 50.221 ;
      RECT 69.677 47.652 69.717 50.221 ;
      RECT 67.193 50.119 69.763 50.175 ;
      RECT 69.69 47.622 69.763 50.175 ;
      RECT 67.239 50.073 69.809 50.129 ;
      RECT 69.736 47.576 69.809 50.129 ;
      RECT 67.285 50.027 69.855 50.083 ;
      RECT 69.782 47.53 69.855 50.083 ;
      RECT 67.331 49.981 69.901 50.037 ;
      RECT 69.828 47.484 69.901 50.037 ;
      RECT 67.377 49.935 69.947 49.991 ;
      RECT 69.874 47.438 69.947 49.991 ;
      RECT 67.423 49.889 69.993 49.945 ;
      RECT 69.92 47.392 69.993 49.945 ;
      RECT 67.469 49.843 70.039 49.899 ;
      RECT 69.966 47.346 70.039 49.899 ;
      RECT 67.515 49.797 70.085 49.853 ;
      RECT 70.012 47.3 70.085 49.853 ;
      RECT 67.561 49.751 70.131 49.807 ;
      RECT 70.058 47.254 70.131 49.807 ;
      RECT 67.607 49.705 70.177 49.761 ;
      RECT 70.104 47.208 70.177 49.761 ;
      RECT 67.653 49.659 70.223 49.715 ;
      RECT 70.15 47.162 70.223 49.715 ;
      RECT 67.699 49.613 70.269 49.669 ;
      RECT 70.196 47.116 70.269 49.669 ;
      RECT 67.745 49.567 70.315 49.623 ;
      RECT 70.242 47.07 70.315 49.623 ;
      RECT 67.791 49.521 70.361 49.577 ;
      RECT 70.288 47.024 70.361 49.577 ;
      RECT 67.837 49.475 70.407 49.531 ;
      RECT 70.334 46.978 70.407 49.531 ;
      RECT 67.883 49.429 70.453 49.485 ;
      RECT 70.38 46.932 70.453 49.485 ;
      RECT 67.929 49.383 70.499 49.439 ;
      RECT 70.426 46.886 70.499 49.439 ;
      RECT 67.975 49.337 70.545 49.393 ;
      RECT 70.472 46.84 70.545 49.393 ;
      RECT 68.021 49.291 70.591 49.347 ;
      RECT 70.518 46.794 70.591 49.347 ;
      RECT 68.067 49.245 70.637 49.301 ;
      RECT 70.564 46.748 70.637 49.301 ;
      RECT 68.113 49.199 70.683 49.255 ;
      RECT 70.61 46.702 70.683 49.255 ;
      RECT 68.159 49.153 70.729 49.209 ;
      RECT 70.656 46.656 70.729 49.209 ;
      RECT 68.205 49.107 70.775 49.163 ;
      RECT 70.702 46.61 70.775 49.163 ;
      RECT 68.251 49.061 70.821 49.117 ;
      RECT 70.748 46.564 70.821 49.117 ;
      RECT 68.297 49.015 70.867 49.071 ;
      RECT 70.794 46.518 70.867 49.071 ;
      RECT 68.343 48.969 70.913 49.025 ;
      RECT 70.84 46.472 70.913 49.025 ;
      RECT 68.389 48.923 70.959 48.979 ;
      RECT 70.886 46.426 70.959 48.979 ;
      RECT 68.435 48.877 71.005 48.933 ;
      RECT 70.932 46.38 71.005 48.933 ;
      RECT 68.481 48.831 71.051 48.887 ;
      RECT 70.978 46.334 71.051 48.887 ;
      RECT 68.527 48.785 71.097 48.841 ;
      RECT 71.024 46.288 71.097 48.841 ;
      RECT 68.573 48.739 71.143 48.795 ;
      RECT 71.07 46.242 71.143 48.795 ;
      RECT 68.619 48.693 71.189 48.749 ;
      RECT 71.116 46.196 71.189 48.749 ;
      RECT 68.665 48.647 71.235 48.703 ;
      RECT 71.162 46.15 71.235 48.703 ;
      RECT 68.711 48.601 71.281 48.657 ;
      RECT 71.208 46.104 71.281 48.657 ;
      RECT 68.757 48.555 71.327 48.611 ;
      RECT 71.254 46.058 71.327 48.611 ;
      RECT 68.803 48.509 71.373 48.565 ;
      RECT 71.3 46.012 71.373 48.565 ;
      RECT 68.849 48.463 71.419 48.519 ;
      RECT 71.346 45.966 71.419 48.519 ;
      RECT 68.895 48.417 71.465 48.473 ;
      RECT 71.392 45.92 71.465 48.473 ;
      RECT 68.941 48.371 71.511 48.427 ;
      RECT 71.438 45.874 71.511 48.427 ;
      RECT 68.987 48.325 71.557 48.381 ;
      RECT 71.484 45.828 71.557 48.381 ;
      RECT 69.033 48.279 71.603 48.335 ;
      RECT 71.53 45.782 71.603 48.335 ;
      RECT 69.079 48.233 71.649 48.289 ;
      RECT 71.576 45.736 71.649 48.289 ;
      RECT 69.125 48.187 71.695 48.243 ;
      RECT 71.622 45.69 71.695 48.243 ;
      RECT 69.171 48.141 71.741 48.197 ;
      RECT 71.668 45.644 71.741 48.197 ;
      RECT 69.217 48.095 71.787 48.151 ;
      RECT 71.714 45.598 71.787 48.151 ;
      RECT 69.263 48.049 71.833 48.105 ;
      RECT 71.76 45.552 71.833 48.105 ;
      RECT 69.309 48.003 71.879 48.059 ;
      RECT 71.806 45.506 71.879 48.059 ;
      RECT 69.355 47.957 71.925 48.013 ;
      RECT 71.852 45.46 71.925 48.013 ;
      RECT 69.401 47.911 71.971 47.967 ;
      RECT 71.898 45.414 71.971 47.967 ;
      RECT 69.447 47.865 72.017 47.921 ;
      RECT 71.944 45.368 72.017 47.921 ;
      RECT 69.493 47.819 72.063 47.875 ;
      RECT 71.99 45.322 72.063 47.875 ;
      RECT 69.539 47.773 72.109 47.829 ;
      RECT 72.036 45.276 72.109 47.829 ;
      RECT 69.585 47.727 72.155 47.783 ;
      RECT 72.082 45.23 72.155 47.783 ;
      RECT 69.631 47.681 72.201 47.737 ;
      RECT 72.128 45.184 72.201 47.737 ;
      RECT 72.174 45.138 72.247 47.691 ;
      RECT 72.22 45.092 72.293 47.645 ;
      RECT 72.266 45.046 72.339 47.599 ;
      RECT 72.312 45 72.385 47.553 ;
      RECT 72.358 44.954 72.431 47.507 ;
      RECT 72.404 44.908 72.477 47.461 ;
      RECT 72.45 44.862 72.523 47.415 ;
      RECT 72.496 44.816 72.569 47.369 ;
      RECT 72.542 44.77 72.615 47.323 ;
      RECT 72.588 44.724 72.661 47.277 ;
      RECT 72.634 44.678 72.707 47.231 ;
      RECT 72.68 44.632 72.753 47.185 ;
      RECT 72.726 44.586 72.799 47.139 ;
      RECT 72.772 44.54 72.845 47.093 ;
      RECT 72.818 44.494 72.891 47.047 ;
      RECT 72.864 44.448 72.937 47.001 ;
      RECT 72.91 44.402 72.983 46.955 ;
      RECT 72.956 44.356 73.029 46.909 ;
      RECT 73.002 44.31 73.075 46.863 ;
      RECT 73.048 44.264 73.121 46.817 ;
      RECT 73.094 44.218 73.167 46.771 ;
      RECT 73.14 44.172 73.213 46.725 ;
      RECT 73.186 44.126 73.259 46.679 ;
      RECT 73.232 44.08 73.305 46.633 ;
      RECT 73.278 44.034 73.351 46.587 ;
      RECT 73.324 43.988 73.397 46.541 ;
      RECT 73.37 43.942 73.443 46.495 ;
      RECT 73.416 43.896 73.489 46.449 ;
      RECT 73.462 43.85 73.535 46.403 ;
      RECT 73.508 43.804 73.581 46.357 ;
      RECT 73.554 43.758 73.627 46.311 ;
      RECT 73.6 43.712 73.673 46.265 ;
      RECT 73.646 43.666 73.719 46.219 ;
      RECT 73.692 43.62 73.765 46.173 ;
      RECT 73.738 43.574 73.811 46.127 ;
      RECT 73.784 43.528 73.857 46.081 ;
      RECT 73.83 43.482 73.903 46.035 ;
      RECT 73.876 43.436 73.949 45.989 ;
      RECT 73.922 43.39 73.995 45.943 ;
      RECT 73.968 43.344 74.041 45.897 ;
      RECT 74.014 43.298 74.087 45.851 ;
      RECT 74.06 43.252 74.133 45.805 ;
      RECT 74.106 43.206 74.179 45.759 ;
      RECT 74.152 43.16 74.225 45.713 ;
      RECT 74.198 43.114 74.271 45.667 ;
      RECT 74.244 43.068 74.317 45.621 ;
      RECT 74.29 43.022 74.363 45.575 ;
      RECT 74.336 42.976 74.409 45.529 ;
      RECT 74.382 42.93 74.455 45.483 ;
      RECT 74.428 42.884 74.501 45.437 ;
      RECT 74.474 42.838 74.547 45.391 ;
      RECT 74.52 42.792 74.593 45.345 ;
      RECT 74.566 42.746 74.639 45.299 ;
      RECT 74.612 42.699 74.685 45.253 ;
      RECT 74.658 42.675 74.731 45.207 ;
      RECT 74.658 42.675 74.777 45.161 ;
      RECT 74.658 42.675 74.823 45.115 ;
      RECT 74.658 42.675 74.869 45.069 ;
      RECT 74.658 42.675 74.915 45.023 ;
      RECT 74.658 42.675 74.961 44.977 ;
      RECT 74.658 42.675 75.007 44.931 ;
      RECT 74.658 42.675 75.053 44.885 ;
      RECT 74.658 42.675 75.099 44.839 ;
      RECT 74.658 42.675 75.145 44.793 ;
      RECT 74.658 42.675 75.191 44.747 ;
      RECT 74.658 42.675 75.237 44.701 ;
      RECT 74.658 42.675 75.283 44.655 ;
      RECT 74.658 42.675 75.329 44.609 ;
      RECT 74.658 42.675 75.375 44.563 ;
      RECT 74.658 42.675 75.421 44.517 ;
      RECT 74.658 42.675 75.467 44.471 ;
      RECT 74.658 42.675 75.513 44.425 ;
      RECT 74.658 42.675 75.559 44.379 ;
      RECT 74.658 42.675 75.605 44.333 ;
      RECT 74.658 42.675 75.651 44.287 ;
      RECT 74.658 42.675 75.697 44.241 ;
      RECT 74.658 42.675 75.743 44.195 ;
      RECT 74.658 42.675 75.789 44.149 ;
      RECT 74.658 42.675 75.835 44.103 ;
      RECT 74.658 42.675 75.881 44.057 ;
      RECT 74.658 42.675 75.927 44.011 ;
      RECT 74.658 42.675 75.973 43.965 ;
      RECT 74.658 42.675 76.019 43.919 ;
      RECT 74.658 42.675 76.065 43.873 ;
      RECT 73.508 43.804 76.09 43.837 ;
      RECT 74.658 42.675 110 43.825 ;
      RECT 56.175 81.387 57.325 110 ;
      RECT 56.175 81.387 57.371 82.562 ;
      RECT 56.175 81.387 57.417 82.516 ;
      RECT 56.175 81.387 57.463 82.47 ;
      RECT 56.175 81.387 57.509 82.424 ;
      RECT 56.175 81.387 57.555 82.378 ;
      RECT 56.175 81.387 57.601 82.332 ;
      RECT 56.175 81.387 57.647 82.286 ;
      RECT 56.175 81.387 57.693 82.24 ;
      RECT 56.175 81.387 57.739 82.194 ;
      RECT 56.175 81.387 57.785 82.148 ;
      RECT 56.175 81.387 57.831 82.102 ;
      RECT 56.175 81.387 57.877 82.056 ;
      RECT 56.175 81.387 57.923 82.01 ;
      RECT 56.175 81.387 57.969 81.964 ;
      RECT 56.175 81.387 58.015 81.918 ;
      RECT 56.175 81.387 58.061 81.872 ;
      RECT 56.175 81.387 58.107 81.826 ;
      RECT 56.175 81.387 58.153 81.78 ;
      RECT 56.175 81.387 58.199 81.734 ;
      RECT 56.175 81.387 58.245 81.688 ;
      RECT 56.175 81.387 58.291 81.642 ;
      RECT 56.175 81.387 58.337 81.596 ;
      RECT 56.175 81.387 58.383 81.55 ;
      RECT 56.175 81.387 58.429 81.504 ;
      RECT 56.175 81.387 58.475 81.458 ;
      RECT 56.221 81.341 58.521 81.412 ;
      RECT 56.267 81.295 58.567 81.366 ;
      RECT 56.313 81.249 58.613 81.32 ;
      RECT 56.359 81.203 58.659 81.274 ;
      RECT 56.405 81.157 58.705 81.228 ;
      RECT 56.451 81.111 58.751 81.182 ;
      RECT 56.497 81.065 58.797 81.136 ;
      RECT 56.543 81.019 58.843 81.09 ;
      RECT 56.589 80.973 58.889 81.044 ;
      RECT 56.635 80.927 58.935 80.998 ;
      RECT 56.681 80.881 58.981 80.952 ;
      RECT 56.727 80.835 59.027 80.906 ;
      RECT 56.773 80.789 59.073 80.86 ;
      RECT 56.819 80.743 59.119 80.814 ;
      RECT 56.865 80.697 59.165 80.768 ;
      RECT 56.911 80.651 59.211 80.722 ;
      RECT 56.957 80.605 59.257 80.676 ;
      RECT 57.003 80.559 59.303 80.63 ;
      RECT 57.049 80.513 59.349 80.584 ;
      RECT 57.095 80.467 59.395 80.538 ;
      RECT 57.141 80.421 59.441 80.492 ;
      RECT 57.187 80.375 59.487 80.446 ;
      RECT 57.233 80.329 59.533 80.4 ;
      RECT 57.279 80.283 59.579 80.354 ;
      RECT 57.325 80.237 59.625 80.308 ;
      RECT 57.371 80.191 59.671 80.262 ;
      RECT 57.417 80.145 59.717 80.216 ;
      RECT 57.463 80.099 59.763 80.17 ;
      RECT 57.509 80.053 59.809 80.124 ;
      RECT 57.555 80.007 59.855 80.078 ;
      RECT 57.601 79.961 59.901 80.032 ;
      RECT 57.647 79.915 59.947 79.986 ;
      RECT 57.693 79.869 59.993 79.94 ;
      RECT 57.739 79.823 60.039 79.894 ;
      RECT 57.785 79.777 60.085 79.848 ;
      RECT 57.831 79.731 60.131 79.802 ;
      RECT 57.877 79.685 60.177 79.756 ;
      RECT 57.923 79.639 60.223 79.71 ;
      RECT 57.969 79.593 60.269 79.664 ;
      RECT 58.015 79.547 60.315 79.618 ;
      RECT 58.061 79.501 60.361 79.572 ;
      RECT 58.107 79.455 60.407 79.526 ;
      RECT 58.153 79.409 60.453 79.48 ;
      RECT 58.199 79.363 60.499 79.434 ;
      RECT 58.245 79.317 60.545 79.388 ;
      RECT 58.291 79.271 60.591 79.342 ;
      RECT 58.337 79.225 60.637 79.296 ;
      RECT 58.383 79.179 60.683 79.25 ;
      RECT 58.429 79.133 60.729 79.204 ;
      RECT 58.475 79.087 60.775 79.158 ;
      RECT 58.521 79.041 60.821 79.112 ;
      RECT 58.567 78.995 60.867 79.066 ;
      RECT 58.613 78.949 60.913 79.02 ;
      RECT 58.659 78.903 60.959 78.974 ;
      RECT 58.705 78.857 61.005 78.928 ;
      RECT 58.751 78.811 61.051 78.882 ;
      RECT 58.797 78.765 61.097 78.836 ;
      RECT 58.843 78.719 61.143 78.79 ;
      RECT 58.889 78.673 61.189 78.744 ;
      RECT 58.935 78.627 61.235 78.698 ;
      RECT 58.981 78.581 61.281 78.652 ;
      RECT 59.027 78.535 61.327 78.606 ;
      RECT 59.073 78.489 61.373 78.56 ;
      RECT 59.119 78.443 61.419 78.514 ;
      RECT 59.165 78.397 61.465 78.468 ;
      RECT 59.211 78.351 61.511 78.422 ;
      RECT 59.257 78.305 61.557 78.376 ;
      RECT 59.303 78.259 61.603 78.33 ;
      RECT 59.349 78.213 61.649 78.284 ;
      RECT 59.395 78.167 61.695 78.238 ;
      RECT 59.441 78.121 61.741 78.192 ;
      RECT 59.487 78.075 61.787 78.146 ;
      RECT 59.533 78.029 61.833 78.1 ;
      RECT 59.579 77.983 61.879 78.054 ;
      RECT 59.625 77.937 61.925 78.008 ;
      RECT 59.671 77.891 61.971 77.962 ;
      RECT 59.717 77.845 62.017 77.916 ;
      RECT 59.763 77.799 62.063 77.87 ;
      RECT 59.809 77.753 62.109 77.824 ;
      RECT 59.855 77.707 62.155 77.778 ;
      RECT 59.901 77.661 62.201 77.732 ;
      RECT 59.947 77.615 62.247 77.686 ;
      RECT 59.993 77.569 62.293 77.64 ;
      RECT 60.039 77.523 62.339 77.594 ;
      RECT 60.085 77.477 62.385 77.548 ;
      RECT 60.131 77.431 62.431 77.502 ;
      RECT 60.177 77.385 62.477 77.456 ;
      RECT 60.223 77.339 62.523 77.41 ;
      RECT 60.269 77.293 62.569 77.364 ;
      RECT 60.315 77.247 62.615 77.318 ;
      RECT 60.361 77.201 62.661 77.272 ;
      RECT 60.407 77.155 62.707 77.226 ;
      RECT 60.453 77.109 62.753 77.18 ;
      RECT 60.499 77.063 62.799 77.134 ;
      RECT 60.545 77.017 62.845 77.088 ;
      RECT 60.591 76.971 62.891 77.042 ;
      RECT 60.637 76.925 62.937 76.996 ;
      RECT 60.683 76.879 62.983 76.95 ;
      RECT 60.729 76.833 63.029 76.904 ;
      RECT 60.775 76.787 63.075 76.858 ;
      RECT 60.821 76.741 63.121 76.812 ;
      RECT 60.867 76.695 63.167 76.766 ;
      RECT 60.913 76.649 63.213 76.72 ;
      RECT 60.959 76.603 63.259 76.674 ;
      RECT 61.005 76.557 63.305 76.628 ;
      RECT 61.005 76.557 63.325 76.595 ;
      RECT 61.051 76.511 63.371 76.562 ;
      RECT 63.305 74.257 63.371 76.562 ;
      RECT 61.097 76.465 63.417 76.516 ;
      RECT 63.351 74.211 63.417 76.516 ;
      RECT 61.143 76.419 63.463 76.47 ;
      RECT 63.397 74.165 63.463 76.47 ;
      RECT 61.189 76.373 63.509 76.424 ;
      RECT 63.443 74.119 63.509 76.424 ;
      RECT 61.235 76.327 63.555 76.378 ;
      RECT 63.489 74.073 63.555 76.378 ;
      RECT 61.281 76.281 63.601 76.332 ;
      RECT 63.535 74.027 63.601 76.332 ;
      RECT 61.327 76.235 63.647 76.286 ;
      RECT 63.581 73.981 63.647 76.286 ;
      RECT 61.373 76.189 63.693 76.24 ;
      RECT 63.627 73.935 63.693 76.24 ;
      RECT 61.419 76.143 63.739 76.194 ;
      RECT 63.673 73.889 63.739 76.194 ;
      RECT 61.465 76.097 63.785 76.148 ;
      RECT 63.719 73.843 63.785 76.148 ;
      RECT 61.511 76.051 63.831 76.102 ;
      RECT 63.765 73.797 63.831 76.102 ;
      RECT 61.557 76.005 63.877 76.056 ;
      RECT 63.811 73.751 63.877 76.056 ;
      RECT 61.603 75.959 63.923 76.01 ;
      RECT 63.857 73.705 63.923 76.01 ;
      RECT 61.649 75.913 63.969 75.964 ;
      RECT 63.903 73.659 63.969 75.964 ;
      RECT 61.695 75.867 64.015 75.918 ;
      RECT 63.949 73.613 64.015 75.918 ;
      RECT 61.741 75.821 64.061 75.872 ;
      RECT 63.995 73.567 64.061 75.872 ;
      RECT 61.787 75.775 64.107 75.826 ;
      RECT 64.041 73.521 64.107 75.826 ;
      RECT 61.833 75.729 64.153 75.78 ;
      RECT 64.087 73.475 64.153 75.78 ;
      RECT 61.879 75.683 64.199 75.734 ;
      RECT 64.133 73.429 64.199 75.734 ;
      RECT 61.925 75.637 64.245 75.688 ;
      RECT 64.179 73.383 64.245 75.688 ;
      RECT 61.971 75.591 64.291 75.642 ;
      RECT 64.225 73.337 64.291 75.642 ;
      RECT 62.017 75.545 64.337 75.596 ;
      RECT 64.271 73.291 64.337 75.596 ;
      RECT 62.063 75.499 64.383 75.55 ;
      RECT 64.317 73.245 64.383 75.55 ;
      RECT 62.109 75.453 64.429 75.504 ;
      RECT 64.363 73.199 64.429 75.504 ;
      RECT 62.155 75.407 64.475 75.458 ;
      RECT 64.409 73.153 64.475 75.458 ;
      RECT 62.201 75.361 64.521 75.412 ;
      RECT 64.455 73.107 64.521 75.412 ;
      RECT 62.247 75.315 64.567 75.366 ;
      RECT 64.501 73.061 64.567 75.366 ;
      RECT 62.293 75.269 64.613 75.32 ;
      RECT 64.547 73.015 64.613 75.32 ;
      RECT 62.339 75.223 64.659 75.274 ;
      RECT 64.593 72.969 64.659 75.274 ;
      RECT 62.385 75.177 64.705 75.228 ;
      RECT 64.639 72.923 64.705 75.228 ;
      RECT 62.431 75.131 64.751 75.182 ;
      RECT 64.685 72.877 64.751 75.182 ;
      RECT 62.477 75.085 64.797 75.136 ;
      RECT 64.731 72.831 64.797 75.136 ;
      RECT 62.523 75.039 64.843 75.09 ;
      RECT 64.777 72.785 64.843 75.09 ;
      RECT 62.569 74.993 64.889 75.044 ;
      RECT 64.823 72.739 64.889 75.044 ;
      RECT 62.615 74.947 64.935 74.998 ;
      RECT 64.869 72.693 64.935 74.998 ;
      RECT 62.661 74.901 64.981 74.952 ;
      RECT 64.915 72.647 64.981 74.952 ;
      RECT 62.707 74.855 65.027 74.906 ;
      RECT 64.961 72.601 65.027 74.906 ;
      RECT 62.753 74.809 65.073 74.86 ;
      RECT 65.007 72.555 65.073 74.86 ;
      RECT 62.799 74.763 65.119 74.814 ;
      RECT 65.053 72.509 65.119 74.814 ;
      RECT 62.845 74.717 65.165 74.768 ;
      RECT 65.099 72.463 65.165 74.768 ;
      RECT 62.891 74.671 65.211 74.722 ;
      RECT 65.145 72.417 65.211 74.722 ;
      RECT 62.937 74.625 65.257 74.676 ;
      RECT 65.191 72.371 65.257 74.676 ;
      RECT 62.983 74.579 65.303 74.63 ;
      RECT 65.237 72.325 65.303 74.63 ;
      RECT 63.029 74.533 65.349 74.584 ;
      RECT 65.283 72.279 65.349 74.584 ;
      RECT 63.075 74.487 65.395 74.538 ;
      RECT 65.329 72.233 65.395 74.538 ;
      RECT 63.121 74.441 65.441 74.492 ;
      RECT 65.375 72.187 65.441 74.492 ;
      RECT 63.167 74.395 65.487 74.446 ;
      RECT 65.421 72.141 65.487 74.446 ;
      RECT 63.213 74.349 65.533 74.4 ;
      RECT 65.467 72.095 65.533 74.4 ;
      RECT 63.259 74.303 65.579 74.354 ;
      RECT 65.513 72.049 65.579 74.354 ;
      RECT 65.559 72.003 65.625 74.308 ;
      RECT 65.605 71.957 65.671 74.262 ;
      RECT 65.651 71.911 65.717 74.216 ;
      RECT 65.697 71.865 65.763 74.17 ;
      RECT 65.743 71.819 65.809 74.124 ;
      RECT 65.789 71.773 65.855 74.078 ;
      RECT 65.835 71.727 65.901 74.032 ;
      RECT 65.881 71.681 65.947 73.986 ;
      RECT 65.927 71.635 65.993 73.94 ;
      RECT 65.973 71.589 66.039 73.894 ;
      RECT 66.019 71.543 66.085 73.848 ;
      RECT 66.065 71.497 66.131 73.802 ;
      RECT 66.111 71.451 66.177 73.756 ;
      RECT 66.157 71.405 66.223 73.71 ;
      RECT 66.203 71.359 66.269 73.664 ;
      RECT 66.249 71.313 66.315 73.618 ;
      RECT 66.295 71.267 66.361 73.572 ;
      RECT 66.341 71.221 66.407 73.526 ;
      RECT 66.387 71.175 66.453 73.48 ;
      RECT 66.433 71.129 66.499 73.434 ;
      RECT 66.479 71.083 66.545 73.388 ;
      RECT 66.525 71.037 66.591 73.342 ;
      RECT 66.571 70.991 66.637 73.296 ;
      RECT 66.617 70.945 66.683 73.25 ;
      RECT 66.663 70.899 66.729 73.204 ;
      RECT 66.709 70.853 66.775 73.158 ;
      RECT 66.755 70.807 66.821 73.112 ;
      RECT 66.801 70.761 66.867 73.066 ;
      RECT 66.847 70.715 66.913 73.02 ;
      RECT 66.893 70.669 66.959 72.974 ;
      RECT 66.939 70.623 67.005 72.928 ;
      RECT 66.985 70.577 67.051 72.882 ;
      RECT 67.031 70.531 67.097 72.836 ;
      RECT 67.077 70.485 67.143 72.79 ;
      RECT 67.123 70.439 67.189 72.744 ;
      RECT 67.169 70.393 67.235 72.698 ;
      RECT 67.215 70.347 67.281 72.652 ;
      RECT 67.261 70.301 67.327 72.606 ;
      RECT 67.307 70.255 67.373 72.56 ;
      RECT 67.353 70.209 67.419 72.514 ;
      RECT 67.399 70.163 67.465 72.468 ;
      RECT 67.445 70.117 67.511 72.422 ;
      RECT 67.491 70.071 67.557 72.376 ;
      RECT 67.537 70.025 67.603 72.33 ;
      RECT 67.583 69.979 67.649 72.284 ;
      RECT 67.629 69.933 67.695 72.238 ;
      RECT 67.675 69.887 67.741 72.192 ;
      RECT 67.721 69.841 67.787 72.146 ;
      RECT 67.767 69.795 67.833 72.1 ;
      RECT 67.813 69.749 67.879 72.054 ;
      RECT 67.859 69.703 67.925 72.008 ;
      RECT 67.905 69.657 67.971 71.962 ;
      RECT 67.951 69.611 68.017 71.916 ;
      RECT 67.997 69.565 68.063 71.87 ;
      RECT 68.043 69.519 68.109 71.824 ;
      RECT 68.089 69.473 68.155 71.778 ;
      RECT 68.135 69.427 68.201 71.732 ;
      RECT 68.181 69.381 68.247 71.686 ;
      RECT 68.227 69.335 68.293 71.64 ;
      RECT 68.273 69.289 68.339 71.594 ;
      RECT 68.319 69.243 68.385 71.548 ;
      RECT 68.365 69.197 68.431 71.502 ;
      RECT 68.411 69.151 68.477 71.456 ;
      RECT 68.457 69.105 68.523 71.41 ;
      RECT 68.503 69.059 68.569 71.364 ;
      RECT 68.549 69.013 68.615 71.318 ;
      RECT 68.595 68.967 68.661 71.272 ;
      RECT 68.641 68.921 68.707 71.226 ;
      RECT 68.687 68.875 68.753 71.18 ;
      RECT 68.733 68.829 68.799 71.134 ;
      RECT 68.779 68.783 68.845 71.088 ;
      RECT 68.825 68.737 68.891 71.042 ;
      RECT 68.871 68.691 68.937 70.996 ;
      RECT 68.917 68.645 68.983 70.95 ;
      RECT 68.963 68.599 69.029 70.904 ;
      RECT 69.009 68.553 69.075 70.858 ;
      RECT 69.055 68.507 69.121 70.812 ;
      RECT 69.101 68.461 69.167 70.766 ;
      RECT 69.147 68.415 69.213 70.72 ;
      RECT 69.193 68.369 69.259 70.674 ;
      RECT 69.239 68.323 69.305 70.628 ;
      RECT 69.285 68.277 69.351 70.582 ;
      RECT 69.331 68.231 69.397 70.536 ;
      RECT 69.377 68.185 69.443 70.49 ;
      RECT 69.423 68.139 69.489 70.444 ;
      RECT 69.469 68.093 69.535 70.398 ;
      RECT 69.515 68.047 69.581 70.352 ;
      RECT 69.561 68.001 69.627 70.306 ;
      RECT 69.607 67.955 69.673 70.26 ;
      RECT 69.653 67.909 69.719 70.214 ;
      RECT 69.699 67.863 69.765 70.168 ;
      RECT 69.745 67.817 69.811 70.122 ;
      RECT 69.791 67.771 69.857 70.076 ;
      RECT 69.837 67.725 69.903 70.03 ;
      RECT 69.883 67.679 69.949 69.984 ;
      RECT 69.929 67.633 69.995 69.938 ;
      RECT 69.975 67.587 70.041 69.892 ;
      RECT 70.021 67.541 70.087 69.846 ;
      RECT 70.067 67.495 70.133 69.8 ;
      RECT 70.113 67.449 70.179 69.754 ;
      RECT 70.159 67.403 70.225 69.708 ;
      RECT 70.205 67.357 70.271 69.662 ;
      RECT 70.251 67.311 70.317 69.616 ;
      RECT 70.297 67.265 70.363 69.57 ;
      RECT 70.343 67.219 70.409 69.524 ;
      RECT 70.389 67.173 70.455 69.478 ;
      RECT 70.435 67.127 70.501 69.432 ;
      RECT 70.481 67.081 70.547 69.386 ;
      RECT 70.527 67.035 70.593 69.34 ;
      RECT 70.573 66.989 70.639 69.294 ;
      RECT 70.619 66.943 70.685 69.248 ;
      RECT 70.665 66.897 70.731 69.202 ;
      RECT 70.711 66.851 70.777 69.156 ;
      RECT 70.757 66.805 70.823 69.11 ;
      RECT 70.803 66.759 70.869 69.064 ;
      RECT 70.849 66.713 70.915 69.018 ;
      RECT 70.895 66.667 70.961 68.972 ;
      RECT 70.941 66.621 71.007 68.926 ;
      RECT 70.987 66.575 71.053 68.88 ;
      RECT 71.033 66.529 71.099 68.834 ;
      RECT 71.079 66.483 71.145 68.788 ;
      RECT 71.125 66.437 71.191 68.742 ;
      RECT 71.171 66.391 71.237 68.696 ;
      RECT 71.217 66.345 71.283 68.65 ;
      RECT 71.263 66.299 71.329 68.604 ;
      RECT 71.309 66.253 71.375 68.558 ;
      RECT 71.355 66.207 71.421 68.512 ;
      RECT 71.401 66.161 71.467 68.466 ;
      RECT 71.447 66.115 71.513 68.42 ;
      RECT 71.493 66.069 71.559 68.374 ;
      RECT 71.539 66.023 71.605 68.328 ;
      RECT 71.585 65.977 71.651 68.282 ;
      RECT 71.631 65.931 71.697 68.236 ;
      RECT 71.677 65.885 71.743 68.19 ;
      RECT 71.723 65.839 71.789 68.144 ;
      RECT 71.769 65.793 71.835 68.098 ;
      RECT 71.815 65.747 71.881 68.052 ;
      RECT 71.861 65.701 71.927 68.006 ;
      RECT 71.907 65.655 71.973 67.96 ;
      RECT 71.953 65.609 72.019 67.914 ;
      RECT 71.999 65.563 72.065 67.868 ;
      RECT 72.045 65.517 72.111 67.822 ;
      RECT 72.091 65.471 72.157 67.776 ;
      RECT 72.137 65.425 72.203 67.73 ;
      RECT 72.183 65.379 72.249 67.684 ;
      RECT 72.229 65.333 72.295 67.638 ;
      RECT 72.275 65.287 72.341 67.592 ;
      RECT 72.321 65.241 72.387 67.546 ;
      RECT 72.367 65.195 72.433 67.5 ;
      RECT 72.413 65.149 72.479 67.454 ;
      RECT 72.459 65.103 72.525 67.408 ;
      RECT 72.505 65.057 72.571 67.362 ;
      RECT 72.551 65.011 72.617 67.316 ;
      RECT 72.597 64.965 72.663 67.27 ;
      RECT 72.643 64.919 72.709 67.224 ;
      RECT 72.689 64.873 72.755 67.178 ;
      RECT 72.735 64.827 72.801 67.132 ;
      RECT 72.781 64.781 72.847 67.086 ;
      RECT 72.827 64.735 72.893 67.04 ;
      RECT 72.873 64.689 72.939 66.994 ;
      RECT 72.919 64.643 72.985 66.948 ;
      RECT 72.965 64.597 73.031 66.902 ;
      RECT 73.011 64.551 73.077 66.856 ;
      RECT 73.057 64.505 73.123 66.81 ;
      RECT 73.103 64.459 73.169 66.764 ;
      RECT 73.149 64.413 73.215 66.718 ;
      RECT 73.195 64.367 73.261 66.672 ;
      RECT 73.241 64.321 73.307 66.626 ;
      RECT 73.287 64.275 73.353 66.58 ;
      RECT 73.333 64.229 73.399 66.534 ;
      RECT 73.379 64.183 73.445 66.488 ;
      RECT 73.425 64.137 73.491 66.442 ;
      RECT 73.471 64.091 73.537 66.396 ;
      RECT 73.517 64.045 73.583 66.35 ;
      RECT 73.563 63.999 73.629 66.304 ;
      RECT 73.609 63.953 73.675 66.258 ;
      RECT 73.655 63.907 73.721 66.212 ;
      RECT 73.701 63.861 73.767 66.166 ;
      RECT 73.747 63.815 73.813 66.12 ;
      RECT 73.793 63.769 73.859 66.074 ;
      RECT 73.839 63.723 73.905 66.028 ;
      RECT 73.885 63.677 73.951 65.982 ;
      RECT 73.931 63.631 73.997 65.936 ;
      RECT 73.977 63.585 74.043 65.89 ;
      RECT 74.023 63.539 74.089 65.844 ;
      RECT 74.069 63.493 74.135 65.798 ;
      RECT 74.115 63.447 74.181 65.752 ;
      RECT 74.161 63.401 74.227 65.706 ;
      RECT 74.207 63.355 74.273 65.66 ;
      RECT 74.253 63.309 74.319 65.614 ;
      RECT 74.299 63.263 74.365 65.568 ;
      RECT 74.345 63.217 74.411 65.522 ;
      RECT 74.391 63.171 74.457 65.476 ;
      RECT 74.437 63.125 74.503 65.43 ;
      RECT 74.483 63.079 74.549 65.384 ;
      RECT 74.529 63.033 74.595 65.338 ;
      RECT 74.575 62.987 74.641 65.292 ;
      RECT 74.621 62.941 74.687 65.246 ;
      RECT 74.667 62.895 74.733 65.2 ;
      RECT 74.713 62.849 74.779 65.154 ;
      RECT 74.759 62.803 74.825 65.108 ;
      RECT 74.805 62.757 74.871 65.062 ;
      RECT 74.851 62.711 74.917 65.016 ;
      RECT 74.897 62.665 74.963 64.97 ;
      RECT 74.943 62.619 75.009 64.924 ;
      RECT 74.989 62.573 75.055 64.878 ;
      RECT 75.035 62.527 75.101 64.832 ;
      RECT 75.081 62.481 75.147 64.786 ;
      RECT 75.127 62.435 75.193 64.74 ;
      RECT 75.173 62.389 75.239 64.694 ;
      RECT 75.219 62.343 75.285 64.648 ;
      RECT 75.265 62.297 75.331 64.602 ;
      RECT 75.311 62.251 75.377 64.556 ;
      RECT 75.357 62.205 75.423 64.51 ;
      RECT 75.403 62.159 75.469 64.464 ;
      RECT 75.449 62.113 75.515 64.418 ;
      RECT 75.495 62.067 75.561 64.372 ;
      RECT 75.541 62.021 75.607 64.326 ;
      RECT 75.587 61.975 75.653 64.28 ;
      RECT 75.633 61.929 75.699 64.234 ;
      RECT 75.679 61.883 75.745 64.188 ;
      RECT 75.725 61.837 75.791 64.142 ;
      RECT 75.771 61.791 75.837 64.096 ;
      RECT 75.817 61.745 75.883 64.05 ;
      RECT 75.863 61.699 75.929 64.004 ;
      RECT 75.909 61.653 75.975 63.958 ;
      RECT 75.955 61.607 76.021 63.912 ;
      RECT 76.001 61.561 76.067 63.866 ;
      RECT 76.047 61.515 76.113 63.82 ;
      RECT 76.093 61.469 76.159 63.774 ;
      RECT 76.139 61.423 76.205 63.728 ;
      RECT 76.185 61.377 76.251 63.682 ;
      RECT 76.231 61.331 76.297 63.636 ;
      RECT 76.277 61.285 76.343 63.59 ;
      RECT 76.323 61.239 76.389 63.544 ;
      RECT 76.369 61.193 76.435 63.498 ;
      RECT 76.415 61.158 76.481 63.452 ;
      RECT 76.44 61.122 76.527 63.406 ;
      RECT 76.486 61.076 76.573 63.36 ;
      RECT 76.532 61.03 76.619 63.314 ;
      RECT 76.578 60.984 76.665 63.268 ;
      RECT 76.624 60.938 76.711 63.222 ;
      RECT 76.67 60.892 76.757 63.176 ;
      RECT 76.716 60.846 76.803 63.13 ;
      RECT 76.762 60.8 76.849 63.084 ;
      RECT 76.808 60.754 76.895 63.038 ;
      RECT 76.854 60.708 76.941 62.992 ;
      RECT 76.9 60.662 76.987 62.946 ;
      RECT 76.946 60.616 77.033 62.9 ;
      RECT 76.992 60.57 77.079 62.854 ;
      RECT 77.038 60.524 77.125 62.808 ;
      RECT 77.084 60.478 77.171 62.762 ;
      RECT 77.13 60.432 77.217 62.716 ;
      RECT 77.176 60.386 77.263 62.67 ;
      RECT 77.222 60.34 77.309 62.624 ;
      RECT 77.268 60.294 77.355 62.578 ;
      RECT 77.314 60.248 77.401 62.532 ;
      RECT 77.36 60.202 77.447 62.486 ;
      RECT 77.406 60.156 77.493 62.44 ;
      RECT 77.452 60.11 77.539 62.394 ;
      RECT 77.498 60.064 77.585 62.348 ;
      RECT 77.544 60.018 77.631 62.302 ;
      RECT 77.59 59.972 77.677 62.256 ;
      RECT 77.636 59.926 77.723 62.21 ;
      RECT 77.682 59.88 77.769 62.164 ;
      RECT 77.728 59.834 77.815 62.118 ;
      RECT 77.774 59.788 77.861 62.072 ;
      RECT 77.82 59.742 77.907 62.026 ;
      RECT 77.866 59.696 77.953 61.98 ;
      RECT 77.912 59.65 77.999 61.934 ;
      RECT 77.958 59.604 78.045 61.888 ;
      RECT 78.004 59.558 78.091 61.842 ;
      RECT 78.05 59.512 78.137 61.796 ;
      RECT 78.096 59.466 78.183 61.75 ;
      RECT 78.142 59.42 78.229 61.704 ;
      RECT 78.188 59.374 78.275 61.658 ;
      RECT 78.234 59.328 78.321 61.612 ;
      RECT 78.28 59.282 78.367 61.566 ;
      RECT 78.326 59.236 78.413 61.52 ;
      RECT 78.372 59.19 78.459 61.474 ;
      RECT 78.418 59.144 78.505 61.428 ;
      RECT 78.464 59.098 78.551 61.382 ;
      RECT 78.51 59.052 78.597 61.336 ;
      RECT 78.556 59.006 78.643 61.29 ;
      RECT 78.602 58.96 78.689 61.244 ;
      RECT 78.648 58.914 78.735 61.198 ;
      RECT 78.694 58.868 78.781 61.152 ;
      RECT 78.74 58.822 78.827 61.106 ;
      RECT 78.786 58.776 78.873 61.06 ;
      RECT 78.832 58.73 78.919 61.014 ;
      RECT 78.878 58.684 78.965 60.968 ;
      RECT 78.924 58.638 79.011 60.922 ;
      RECT 78.97 58.592 79.057 60.876 ;
      RECT 79.016 58.546 79.103 60.83 ;
      RECT 79.062 58.5 79.149 60.784 ;
      RECT 79.108 58.454 79.195 60.738 ;
      RECT 79.154 58.408 79.241 60.692 ;
      RECT 79.2 58.362 79.287 60.646 ;
      RECT 79.246 58.316 79.333 60.6 ;
      RECT 79.292 58.27 79.379 60.554 ;
      RECT 79.338 58.224 79.425 60.508 ;
      RECT 79.384 58.178 79.471 60.462 ;
      RECT 79.43 58.132 79.517 60.416 ;
      RECT 79.476 58.086 79.563 60.37 ;
      RECT 79.522 58.04 79.609 60.324 ;
      RECT 79.568 57.994 79.655 60.278 ;
      RECT 79.614 57.948 79.701 60.232 ;
      RECT 79.66 57.902 79.747 60.186 ;
      RECT 79.706 57.856 79.793 60.14 ;
      RECT 79.752 57.81 79.839 60.094 ;
      RECT 79.798 57.764 79.885 60.048 ;
      RECT 79.844 57.718 79.931 60.002 ;
      RECT 79.89 57.672 79.977 59.956 ;
      RECT 79.936 57.626 80.023 59.91 ;
      RECT 79.982 57.58 80.069 59.864 ;
      RECT 80.028 57.534 80.115 59.818 ;
      RECT 80.074 57.488 80.161 59.772 ;
      RECT 80.12 57.442 80.207 59.726 ;
      RECT 80.166 57.396 80.253 59.68 ;
      RECT 80.212 57.35 80.299 59.634 ;
      RECT 80.258 57.304 80.345 59.588 ;
      RECT 80.304 57.258 80.391 59.542 ;
      RECT 80.35 57.212 80.437 59.496 ;
      RECT 80.396 57.166 80.483 59.45 ;
      RECT 80.442 57.12 80.529 59.404 ;
      RECT 80.488 57.074 80.575 59.358 ;
      RECT 80.534 57.028 80.621 59.312 ;
      RECT 80.58 56.982 80.667 59.266 ;
      RECT 80.626 56.936 80.713 59.22 ;
      RECT 80.672 56.89 80.759 59.174 ;
      RECT 80.718 56.844 80.805 59.128 ;
      RECT 80.764 56.798 80.851 59.082 ;
      RECT 80.81 56.752 80.897 59.036 ;
      RECT 80.856 56.706 80.943 58.99 ;
      RECT 80.902 56.66 80.989 58.944 ;
      RECT 80.948 56.614 81.035 58.898 ;
      RECT 80.994 56.568 81.081 58.852 ;
      RECT 81.04 56.522 81.127 58.806 ;
      RECT 81.086 56.476 81.173 58.76 ;
      RECT 81.132 56.43 81.219 58.714 ;
      RECT 81.178 56.384 81.265 58.668 ;
      RECT 81.224 56.338 81.311 58.622 ;
      RECT 81.27 56.292 81.357 58.576 ;
      RECT 81.316 56.246 81.403 58.53 ;
      RECT 81.362 56.199 81.449 58.484 ;
      RECT 81.408 56.175 81.495 58.438 ;
      RECT 81.408 56.175 81.541 58.392 ;
      RECT 81.408 56.175 81.587 58.346 ;
      RECT 81.408 56.175 81.633 58.3 ;
      RECT 81.408 56.175 81.679 58.254 ;
      RECT 81.408 56.175 81.725 58.208 ;
      RECT 81.408 56.175 81.771 58.162 ;
      RECT 81.408 56.175 81.817 58.116 ;
      RECT 81.408 56.175 81.863 58.07 ;
      RECT 81.408 56.175 81.909 58.024 ;
      RECT 81.408 56.175 81.955 57.978 ;
      RECT 81.408 56.175 82.001 57.932 ;
      RECT 81.408 56.175 82.047 57.886 ;
      RECT 81.408 56.175 82.093 57.84 ;
      RECT 81.408 56.175 82.139 57.794 ;
      RECT 81.408 56.175 82.185 57.748 ;
      RECT 81.408 56.175 82.231 57.702 ;
      RECT 81.408 56.175 82.277 57.656 ;
      RECT 81.408 56.175 82.323 57.61 ;
      RECT 81.408 56.175 82.369 57.564 ;
      RECT 81.408 56.175 82.415 57.518 ;
      RECT 81.408 56.175 82.461 57.472 ;
      RECT 81.408 56.175 82.507 57.426 ;
      RECT 81.408 56.175 82.553 57.38 ;
      RECT 80.258 57.304 82.585 57.341 ;
      RECT 81.408 56.175 110 57.325 ;
      RECT 63.675 85.392 68.325 110 ;
      RECT 63.675 85.392 68.371 88.167 ;
      RECT 63.675 85.392 68.417 88.121 ;
      RECT 63.675 85.392 68.463 88.075 ;
      RECT 63.675 85.392 68.509 88.029 ;
      RECT 63.675 85.392 68.555 87.983 ;
      RECT 63.675 85.392 68.601 87.937 ;
      RECT 63.675 85.392 68.647 87.891 ;
      RECT 63.675 85.392 68.693 87.845 ;
      RECT 63.675 85.392 68.739 87.799 ;
      RECT 63.675 85.392 68.785 87.753 ;
      RECT 63.675 85.392 68.831 87.707 ;
      RECT 63.675 85.392 68.877 87.661 ;
      RECT 63.675 85.392 68.923 87.615 ;
      RECT 63.675 85.392 68.969 87.569 ;
      RECT 63.675 85.392 69.015 87.523 ;
      RECT 63.675 85.392 69.061 87.477 ;
      RECT 63.675 85.392 69.107 87.431 ;
      RECT 63.675 85.392 69.153 87.385 ;
      RECT 63.675 85.392 69.199 87.339 ;
      RECT 63.675 85.392 69.245 87.293 ;
      RECT 63.675 85.392 69.291 87.247 ;
      RECT 63.675 85.392 69.337 87.201 ;
      RECT 63.675 85.392 69.383 87.155 ;
      RECT 63.675 85.392 69.429 87.109 ;
      RECT 63.675 85.392 69.475 87.063 ;
      RECT 63.675 85.392 69.521 87.017 ;
      RECT 63.675 85.392 69.567 86.971 ;
      RECT 63.675 85.392 69.613 86.925 ;
      RECT 63.675 85.392 69.659 86.879 ;
      RECT 63.675 85.392 69.705 86.833 ;
      RECT 63.675 85.392 69.751 86.787 ;
      RECT 63.675 85.392 69.797 86.741 ;
      RECT 63.675 85.392 69.843 86.695 ;
      RECT 63.675 85.392 69.889 86.649 ;
      RECT 63.675 85.392 69.935 86.603 ;
      RECT 63.675 85.392 69.981 86.557 ;
      RECT 63.675 85.392 70.027 86.511 ;
      RECT 63.675 85.392 70.073 86.465 ;
      RECT 63.675 85.392 70.119 86.419 ;
      RECT 63.675 85.392 70.165 86.373 ;
      RECT 63.675 85.392 70.211 86.327 ;
      RECT 63.675 85.392 70.257 86.281 ;
      RECT 63.675 85.392 70.303 86.235 ;
      RECT 63.675 85.392 70.349 86.189 ;
      RECT 63.675 85.392 70.395 86.143 ;
      RECT 63.675 85.392 70.441 86.097 ;
      RECT 63.675 85.392 70.487 86.051 ;
      RECT 63.675 85.392 70.533 86.005 ;
      RECT 63.675 85.392 70.579 85.959 ;
      RECT 63.675 85.392 70.625 85.913 ;
      RECT 63.675 85.392 70.671 85.867 ;
      RECT 63.675 85.392 70.717 85.821 ;
      RECT 63.675 85.392 70.763 85.775 ;
      RECT 63.675 85.392 70.809 85.729 ;
      RECT 63.675 85.392 70.855 85.683 ;
      RECT 63.675 85.392 70.901 85.637 ;
      RECT 63.675 85.392 70.947 85.591 ;
      RECT 63.675 85.392 70.993 85.545 ;
      RECT 63.675 85.392 71.039 85.499 ;
      RECT 63.721 85.346 71.131 85.407 ;
      RECT 71.081 77.986 71.131 85.407 ;
      RECT 63.767 85.3 71.177 85.361 ;
      RECT 71.127 77.94 71.177 85.361 ;
      RECT 63.813 85.254 71.223 85.315 ;
      RECT 71.173 77.894 71.223 85.315 ;
      RECT 63.859 85.208 71.269 85.269 ;
      RECT 71.219 77.848 71.269 85.269 ;
      RECT 63.905 85.162 71.315 85.223 ;
      RECT 71.265 77.802 71.315 85.223 ;
      RECT 63.951 85.116 71.361 85.177 ;
      RECT 71.311 77.756 71.361 85.177 ;
      RECT 63.997 85.07 71.407 85.131 ;
      RECT 71.357 77.71 71.407 85.131 ;
      RECT 64.043 85.024 71.453 85.085 ;
      RECT 71.403 77.664 71.453 85.085 ;
      RECT 64.089 84.978 71.499 85.039 ;
      RECT 71.449 77.618 71.499 85.039 ;
      RECT 64.135 84.932 71.545 84.993 ;
      RECT 71.495 77.572 71.545 84.993 ;
      RECT 64.181 84.886 71.591 84.947 ;
      RECT 71.541 77.526 71.591 84.947 ;
      RECT 64.227 84.84 71.637 84.901 ;
      RECT 71.587 77.48 71.637 84.901 ;
      RECT 64.273 84.794 71.683 84.855 ;
      RECT 71.633 77.434 71.683 84.855 ;
      RECT 64.319 84.748 71.729 84.809 ;
      RECT 71.679 77.388 71.729 84.809 ;
      RECT 64.365 84.702 71.775 84.763 ;
      RECT 71.725 77.342 71.775 84.763 ;
      RECT 64.411 84.656 71.821 84.717 ;
      RECT 71.771 77.296 71.821 84.717 ;
      RECT 64.457 84.61 71.867 84.671 ;
      RECT 71.817 77.25 71.867 84.671 ;
      RECT 64.503 84.564 71.913 84.625 ;
      RECT 71.863 77.204 71.913 84.625 ;
      RECT 64.549 84.518 71.959 84.579 ;
      RECT 71.909 77.158 71.959 84.579 ;
      RECT 64.595 84.472 72.005 84.533 ;
      RECT 71.955 77.112 72.005 84.533 ;
      RECT 64.641 84.426 72.051 84.487 ;
      RECT 72.001 77.066 72.051 84.487 ;
      RECT 64.687 84.38 72.097 84.441 ;
      RECT 72.047 77.02 72.097 84.441 ;
      RECT 64.733 84.334 72.143 84.395 ;
      RECT 72.093 76.974 72.143 84.395 ;
      RECT 64.779 84.288 72.189 84.349 ;
      RECT 72.139 76.928 72.189 84.349 ;
      RECT 64.825 84.242 72.235 84.303 ;
      RECT 72.185 76.882 72.235 84.303 ;
      RECT 64.871 84.196 72.281 84.257 ;
      RECT 72.231 76.836 72.281 84.257 ;
      RECT 64.917 84.15 72.327 84.211 ;
      RECT 72.277 76.79 72.327 84.211 ;
      RECT 64.963 84.104 72.373 84.165 ;
      RECT 72.323 76.744 72.373 84.165 ;
      RECT 65.009 84.058 72.419 84.119 ;
      RECT 72.369 76.698 72.419 84.119 ;
      RECT 65.055 84.012 72.465 84.073 ;
      RECT 72.415 76.652 72.465 84.073 ;
      RECT 65.101 83.966 72.511 84.027 ;
      RECT 72.461 76.606 72.511 84.027 ;
      RECT 65.147 83.92 72.557 83.981 ;
      RECT 72.507 76.56 72.557 83.981 ;
      RECT 65.193 83.874 72.603 83.935 ;
      RECT 72.553 76.514 72.603 83.935 ;
      RECT 65.239 83.828 72.649 83.889 ;
      RECT 72.599 76.468 72.649 83.889 ;
      RECT 65.285 83.782 72.695 83.843 ;
      RECT 72.645 76.422 72.695 83.843 ;
      RECT 65.331 83.736 72.741 83.797 ;
      RECT 72.691 76.376 72.741 83.797 ;
      RECT 65.377 83.69 72.787 83.751 ;
      RECT 72.737 76.33 72.787 83.751 ;
      RECT 65.423 83.644 72.833 83.705 ;
      RECT 72.783 76.284 72.833 83.705 ;
      RECT 65.469 83.598 72.879 83.659 ;
      RECT 72.829 76.238 72.879 83.659 ;
      RECT 65.515 83.552 72.925 83.613 ;
      RECT 72.875 76.192 72.925 83.613 ;
      RECT 65.561 83.506 72.971 83.567 ;
      RECT 72.921 76.146 72.971 83.567 ;
      RECT 65.607 83.46 73.017 83.521 ;
      RECT 72.967 76.1 73.017 83.521 ;
      RECT 65.653 83.414 73.063 83.475 ;
      RECT 73.013 76.054 73.063 83.475 ;
      RECT 65.699 83.368 73.109 83.429 ;
      RECT 73.059 76.008 73.109 83.429 ;
      RECT 65.745 83.322 73.155 83.383 ;
      RECT 73.105 75.962 73.155 83.383 ;
      RECT 65.791 83.276 73.201 83.337 ;
      RECT 73.151 75.916 73.201 83.337 ;
      RECT 65.837 83.23 73.247 83.291 ;
      RECT 73.197 75.87 73.247 83.291 ;
      RECT 65.883 83.184 73.293 83.245 ;
      RECT 73.243 75.824 73.293 83.245 ;
      RECT 65.929 83.138 73.339 83.199 ;
      RECT 73.289 75.778 73.339 83.199 ;
      RECT 65.975 83.092 73.385 83.153 ;
      RECT 73.335 75.732 73.385 83.153 ;
      RECT 66.021 83.046 73.431 83.107 ;
      RECT 73.381 75.686 73.431 83.107 ;
      RECT 66.067 83 73.477 83.061 ;
      RECT 73.427 75.64 73.477 83.061 ;
      RECT 66.113 82.954 73.523 83.015 ;
      RECT 73.473 75.594 73.523 83.015 ;
      RECT 66.159 82.908 73.569 82.969 ;
      RECT 73.519 75.548 73.569 82.969 ;
      RECT 66.205 82.862 73.615 82.923 ;
      RECT 73.565 75.502 73.615 82.923 ;
      RECT 66.251 82.816 73.661 82.877 ;
      RECT 73.611 75.456 73.661 82.877 ;
      RECT 66.297 82.77 73.707 82.831 ;
      RECT 73.657 75.41 73.707 82.831 ;
      RECT 66.343 82.724 73.753 82.785 ;
      RECT 73.703 75.364 73.753 82.785 ;
      RECT 66.389 82.678 73.799 82.739 ;
      RECT 73.749 75.318 73.799 82.739 ;
      RECT 66.435 82.632 73.845 82.693 ;
      RECT 73.795 75.272 73.845 82.693 ;
      RECT 66.481 82.586 73.891 82.647 ;
      RECT 73.841 75.226 73.891 82.647 ;
      RECT 66.527 82.54 73.937 82.601 ;
      RECT 73.887 75.18 73.937 82.601 ;
      RECT 66.573 82.494 73.983 82.555 ;
      RECT 73.933 75.134 73.983 82.555 ;
      RECT 66.619 82.448 74.029 82.509 ;
      RECT 73.979 75.088 74.029 82.509 ;
      RECT 66.665 82.402 74.075 82.463 ;
      RECT 74.025 75.042 74.075 82.463 ;
      RECT 66.711 82.356 74.121 82.417 ;
      RECT 74.071 74.996 74.121 82.417 ;
      RECT 66.757 82.31 74.167 82.371 ;
      RECT 74.117 74.95 74.167 82.371 ;
      RECT 66.803 82.264 74.213 82.325 ;
      RECT 74.163 74.904 74.213 82.325 ;
      RECT 66.849 82.218 74.259 82.279 ;
      RECT 74.209 74.858 74.259 82.279 ;
      RECT 66.895 82.172 74.305 82.233 ;
      RECT 74.255 74.812 74.305 82.233 ;
      RECT 66.941 82.126 74.351 82.187 ;
      RECT 74.301 74.766 74.351 82.187 ;
      RECT 66.987 82.08 74.397 82.141 ;
      RECT 74.347 74.72 74.397 82.141 ;
      RECT 67.033 82.034 74.443 82.095 ;
      RECT 74.393 74.674 74.443 82.095 ;
      RECT 67.079 81.988 74.489 82.049 ;
      RECT 74.439 74.628 74.489 82.049 ;
      RECT 67.125 81.942 74.535 82.003 ;
      RECT 74.485 74.582 74.535 82.003 ;
      RECT 67.171 81.896 74.581 81.957 ;
      RECT 74.531 74.536 74.581 81.957 ;
      RECT 67.217 81.85 74.627 81.911 ;
      RECT 74.577 74.49 74.627 81.911 ;
      RECT 67.263 81.804 74.673 81.865 ;
      RECT 74.623 74.444 74.673 81.865 ;
      RECT 67.309 81.758 74.719 81.819 ;
      RECT 74.669 74.398 74.719 81.819 ;
      RECT 67.355 81.712 74.765 81.773 ;
      RECT 74.715 74.352 74.765 81.773 ;
      RECT 67.401 81.666 74.811 81.727 ;
      RECT 74.761 74.306 74.811 81.727 ;
      RECT 67.447 81.62 74.857 81.681 ;
      RECT 74.807 74.26 74.857 81.681 ;
      RECT 67.493 81.574 74.903 81.635 ;
      RECT 74.853 74.214 74.903 81.635 ;
      RECT 67.539 81.528 74.949 81.589 ;
      RECT 74.899 74.168 74.949 81.589 ;
      RECT 67.585 81.482 74.995 81.543 ;
      RECT 74.945 74.122 74.995 81.543 ;
      RECT 67.631 81.436 75.041 81.497 ;
      RECT 74.991 74.076 75.041 81.497 ;
      RECT 67.677 81.39 75.087 81.451 ;
      RECT 75.037 74.03 75.087 81.451 ;
      RECT 67.723 81.344 75.133 81.405 ;
      RECT 75.083 73.984 75.133 81.405 ;
      RECT 67.769 81.298 75.179 81.359 ;
      RECT 75.129 73.938 75.179 81.359 ;
      RECT 67.815 81.252 75.225 81.313 ;
      RECT 75.175 73.892 75.225 81.313 ;
      RECT 67.861 81.206 75.271 81.267 ;
      RECT 75.221 73.846 75.271 81.267 ;
      RECT 67.907 81.16 75.317 81.221 ;
      RECT 75.267 73.8 75.317 81.221 ;
      RECT 67.953 81.114 75.363 81.175 ;
      RECT 75.313 73.754 75.363 81.175 ;
      RECT 67.999 81.068 75.409 81.129 ;
      RECT 75.359 73.708 75.409 81.129 ;
      RECT 68.045 81.022 75.455 81.083 ;
      RECT 75.405 73.662 75.455 81.083 ;
      RECT 68.091 80.976 75.501 81.037 ;
      RECT 75.451 73.616 75.501 81.037 ;
      RECT 68.137 80.93 75.547 80.991 ;
      RECT 75.497 73.57 75.547 80.991 ;
      RECT 68.183 80.884 75.593 80.945 ;
      RECT 75.543 73.524 75.593 80.945 ;
      RECT 68.229 80.838 75.639 80.899 ;
      RECT 75.589 73.478 75.639 80.899 ;
      RECT 68.275 80.792 75.685 80.853 ;
      RECT 75.635 73.432 75.685 80.853 ;
      RECT 68.321 80.746 75.731 80.807 ;
      RECT 75.681 73.386 75.731 80.807 ;
      RECT 68.367 80.7 75.777 80.761 ;
      RECT 75.727 73.34 75.777 80.761 ;
      RECT 68.413 80.654 75.823 80.715 ;
      RECT 75.773 73.294 75.823 80.715 ;
      RECT 68.459 80.608 75.869 80.669 ;
      RECT 75.819 73.248 75.869 80.669 ;
      RECT 68.505 80.562 75.915 80.623 ;
      RECT 75.865 73.202 75.915 80.623 ;
      RECT 68.551 80.516 75.961 80.577 ;
      RECT 75.911 73.156 75.961 80.577 ;
      RECT 68.597 80.47 76.007 80.531 ;
      RECT 75.957 73.11 76.007 80.531 ;
      RECT 68.643 80.424 76.053 80.485 ;
      RECT 76.003 73.064 76.053 80.485 ;
      RECT 68.689 80.378 76.099 80.439 ;
      RECT 76.049 73.018 76.099 80.439 ;
      RECT 68.735 80.332 76.145 80.393 ;
      RECT 76.095 72.972 76.145 80.393 ;
      RECT 68.781 80.286 76.191 80.347 ;
      RECT 76.141 72.926 76.191 80.347 ;
      RECT 68.827 80.24 76.237 80.301 ;
      RECT 76.187 72.88 76.237 80.301 ;
      RECT 68.873 80.194 76.283 80.255 ;
      RECT 76.233 72.834 76.283 80.255 ;
      RECT 68.919 80.148 76.329 80.209 ;
      RECT 76.279 72.788 76.329 80.209 ;
      RECT 68.965 80.102 76.375 80.163 ;
      RECT 76.325 72.742 76.375 80.163 ;
      RECT 69.011 80.056 76.421 80.117 ;
      RECT 76.371 72.696 76.421 80.117 ;
      RECT 69.057 80.01 76.467 80.071 ;
      RECT 76.417 72.65 76.467 80.071 ;
      RECT 69.103 79.964 76.513 80.025 ;
      RECT 76.463 72.604 76.513 80.025 ;
      RECT 69.149 79.918 76.559 79.979 ;
      RECT 76.509 72.558 76.559 79.979 ;
      RECT 69.195 79.872 76.605 79.933 ;
      RECT 76.555 72.512 76.605 79.933 ;
      RECT 69.241 79.826 76.651 79.887 ;
      RECT 76.601 72.466 76.651 79.887 ;
      RECT 69.287 79.78 76.697 79.841 ;
      RECT 76.647 72.42 76.697 79.841 ;
      RECT 69.333 79.734 76.743 79.795 ;
      RECT 76.693 72.374 76.743 79.795 ;
      RECT 69.379 79.688 76.789 79.749 ;
      RECT 76.739 72.328 76.789 79.749 ;
      RECT 69.425 79.642 76.825 79.708 ;
      RECT 71.035 78.032 71.085 85.453 ;
      RECT 69.471 79.596 76.871 79.667 ;
      RECT 76.785 72.282 76.871 79.667 ;
      RECT 69.517 79.55 76.917 79.621 ;
      RECT 76.831 72.236 76.917 79.621 ;
      RECT 69.563 79.504 76.963 79.575 ;
      RECT 76.877 72.19 76.963 79.575 ;
      RECT 69.609 79.458 77.009 79.529 ;
      RECT 76.923 72.144 77.009 79.529 ;
      RECT 69.655 79.412 77.055 79.483 ;
      RECT 76.969 72.098 77.055 79.483 ;
      RECT 69.701 79.366 77.101 79.437 ;
      RECT 77.015 72.052 77.101 79.437 ;
      RECT 69.747 79.32 77.147 79.391 ;
      RECT 77.061 72.006 77.147 79.391 ;
      RECT 69.793 79.274 77.193 79.345 ;
      RECT 77.107 71.96 77.193 79.345 ;
      RECT 69.839 79.228 77.239 79.299 ;
      RECT 77.153 71.914 77.239 79.299 ;
      RECT 69.885 79.182 77.285 79.253 ;
      RECT 77.199 71.868 77.285 79.253 ;
      RECT 69.931 79.136 77.331 79.207 ;
      RECT 77.245 71.822 77.331 79.207 ;
      RECT 69.977 79.09 77.377 79.161 ;
      RECT 77.291 71.776 77.377 79.161 ;
      RECT 70.023 79.044 77.423 79.115 ;
      RECT 77.337 71.73 77.423 79.115 ;
      RECT 70.069 78.998 77.469 79.069 ;
      RECT 77.383 71.684 77.469 79.069 ;
      RECT 70.115 78.952 77.515 79.023 ;
      RECT 77.429 71.638 77.515 79.023 ;
      RECT 70.161 78.906 77.561 78.977 ;
      RECT 77.475 71.592 77.561 78.977 ;
      RECT 70.207 78.86 77.607 78.931 ;
      RECT 77.521 71.546 77.607 78.931 ;
      RECT 70.253 78.814 77.653 78.885 ;
      RECT 77.567 71.5 77.653 78.885 ;
      RECT 70.299 78.768 77.699 78.839 ;
      RECT 77.613 71.454 77.699 78.839 ;
      RECT 70.345 78.722 77.745 78.793 ;
      RECT 77.659 71.408 77.745 78.793 ;
      RECT 70.391 78.676 77.791 78.747 ;
      RECT 77.705 71.362 77.791 78.747 ;
      RECT 70.437 78.63 77.837 78.701 ;
      RECT 77.751 71.316 77.837 78.701 ;
      RECT 70.483 78.584 77.883 78.655 ;
      RECT 77.797 71.27 77.883 78.655 ;
      RECT 70.529 78.538 77.929 78.609 ;
      RECT 77.843 71.224 77.929 78.609 ;
      RECT 70.575 78.492 77.975 78.563 ;
      RECT 77.889 71.178 77.975 78.563 ;
      RECT 70.621 78.446 78.021 78.517 ;
      RECT 77.935 71.132 78.021 78.517 ;
      RECT 70.667 78.4 78.067 78.471 ;
      RECT 77.981 71.086 78.067 78.471 ;
      RECT 70.713 78.354 78.113 78.425 ;
      RECT 78.027 71.04 78.113 78.425 ;
      RECT 70.759 78.308 78.159 78.379 ;
      RECT 78.073 70.994 78.159 78.379 ;
      RECT 70.805 78.262 78.205 78.333 ;
      RECT 78.119 70.948 78.205 78.333 ;
      RECT 70.851 78.216 78.251 78.287 ;
      RECT 78.165 70.902 78.251 78.287 ;
      RECT 70.897 78.17 78.297 78.241 ;
      RECT 78.211 70.856 78.297 78.241 ;
      RECT 70.943 78.124 78.343 78.195 ;
      RECT 78.257 70.81 78.343 78.195 ;
      RECT 70.989 78.078 78.389 78.149 ;
      RECT 78.303 70.764 78.389 78.149 ;
      RECT 78.349 70.718 78.435 78.103 ;
      RECT 78.395 70.672 78.481 78.057 ;
      RECT 78.441 70.626 78.527 78.011 ;
      RECT 78.487 70.58 78.573 77.965 ;
      RECT 78.533 70.534 78.619 77.919 ;
      RECT 78.579 70.488 78.665 77.873 ;
      RECT 78.625 70.442 78.711 77.827 ;
      RECT 78.671 70.396 78.757 77.781 ;
      RECT 78.717 70.35 78.803 77.735 ;
      RECT 78.763 70.304 78.849 77.689 ;
      RECT 78.809 70.258 78.895 77.643 ;
      RECT 78.855 70.212 78.941 77.597 ;
      RECT 78.901 70.166 78.987 77.551 ;
      RECT 78.947 70.12 79.033 77.505 ;
      RECT 78.993 70.074 79.079 77.459 ;
      RECT 79.039 70.028 79.125 77.413 ;
      RECT 79.085 69.982 79.171 77.367 ;
      RECT 79.131 69.936 79.217 77.321 ;
      RECT 79.177 69.89 79.263 77.275 ;
      RECT 79.223 69.844 79.309 77.229 ;
      RECT 79.269 69.798 79.355 77.183 ;
      RECT 79.315 69.752 79.401 77.137 ;
      RECT 79.361 69.706 79.447 77.091 ;
      RECT 79.407 69.66 79.493 77.045 ;
      RECT 79.453 69.614 79.539 76.999 ;
      RECT 79.499 69.568 79.585 76.953 ;
      RECT 79.545 69.522 79.631 76.907 ;
      RECT 79.591 69.476 79.677 76.861 ;
      RECT 79.637 69.43 79.723 76.815 ;
      RECT 79.683 69.384 79.769 76.769 ;
      RECT 79.729 69.338 79.815 76.723 ;
      RECT 79.775 69.292 79.861 76.677 ;
      RECT 79.821 69.246 79.907 76.631 ;
      RECT 79.867 69.2 79.953 76.585 ;
      RECT 79.913 69.154 79.999 76.539 ;
      RECT 79.959 69.108 80.045 76.493 ;
      RECT 80.005 69.062 80.091 76.447 ;
      RECT 80.051 69.016 80.137 76.401 ;
      RECT 80.097 68.97 80.183 76.355 ;
      RECT 80.143 68.924 80.229 76.309 ;
      RECT 80.189 68.878 80.275 76.263 ;
      RECT 80.235 68.832 80.321 76.217 ;
      RECT 80.281 68.786 80.367 76.171 ;
      RECT 80.327 68.74 80.413 76.125 ;
      RECT 80.373 68.694 80.459 76.079 ;
      RECT 80.419 68.648 80.505 76.033 ;
      RECT 80.465 68.602 80.551 75.987 ;
      RECT 80.511 68.556 80.597 75.941 ;
      RECT 80.557 68.51 80.643 75.895 ;
      RECT 80.603 68.464 80.689 75.849 ;
      RECT 80.649 68.418 80.735 75.803 ;
      RECT 80.695 68.372 80.781 75.757 ;
      RECT 80.741 68.326 80.827 75.711 ;
      RECT 80.787 68.28 80.873 75.665 ;
      RECT 80.833 68.234 80.919 75.619 ;
      RECT 80.879 68.188 80.965 75.573 ;
      RECT 80.925 68.142 81.011 75.527 ;
      RECT 80.971 68.096 81.057 75.481 ;
      RECT 81.017 68.05 81.103 75.435 ;
      RECT 81.063 68.004 81.149 75.389 ;
      RECT 81.109 67.958 81.195 75.343 ;
      RECT 81.155 67.912 81.241 75.297 ;
      RECT 81.201 67.866 81.287 75.251 ;
      RECT 81.247 67.82 81.333 75.205 ;
      RECT 81.293 67.774 81.379 75.159 ;
      RECT 81.339 67.728 81.425 75.113 ;
      RECT 81.385 67.682 81.471 75.067 ;
      RECT 81.431 67.636 81.517 75.021 ;
      RECT 81.477 67.59 81.563 74.975 ;
      RECT 81.523 67.544 81.609 74.929 ;
      RECT 81.569 67.498 81.655 74.883 ;
      RECT 81.615 67.452 81.701 74.837 ;
      RECT 81.661 67.406 81.747 74.791 ;
      RECT 81.707 67.36 81.793 74.745 ;
      RECT 81.753 67.314 81.839 74.699 ;
      RECT 81.799 67.268 81.885 74.653 ;
      RECT 81.845 67.222 81.931 74.607 ;
      RECT 81.891 67.176 81.977 74.561 ;
      RECT 81.937 67.13 82.023 74.515 ;
      RECT 81.983 67.084 82.069 74.469 ;
      RECT 82.029 67.038 82.115 74.423 ;
      RECT 82.075 66.992 82.161 74.377 ;
      RECT 82.121 66.946 82.207 74.331 ;
      RECT 82.167 66.9 82.253 74.285 ;
      RECT 82.213 66.854 82.299 74.239 ;
      RECT 82.259 66.808 82.345 74.193 ;
      RECT 82.305 66.762 82.391 74.147 ;
      RECT 82.351 66.716 82.437 74.101 ;
      RECT 82.397 66.67 82.483 74.055 ;
      RECT 82.443 66.624 82.529 74.009 ;
      RECT 82.489 66.578 82.575 73.963 ;
      RECT 82.535 66.532 82.621 73.917 ;
      RECT 82.581 66.486 82.667 73.871 ;
      RECT 82.627 66.44 82.713 73.825 ;
      RECT 82.673 66.394 82.759 73.779 ;
      RECT 82.719 66.348 82.805 73.733 ;
      RECT 82.765 66.302 82.851 73.687 ;
      RECT 82.811 66.256 82.897 73.641 ;
      RECT 82.903 66.171 82.943 73.595 ;
      RECT 82.935 66.132 82.989 73.549 ;
      RECT 82.981 66.086 83.035 73.503 ;
      RECT 83.027 66.04 83.081 73.457 ;
      RECT 83.073 65.994 83.127 73.411 ;
      RECT 83.119 65.948 83.173 73.365 ;
      RECT 83.165 65.902 83.219 73.319 ;
      RECT 83.211 65.856 83.265 73.273 ;
      RECT 83.257 65.81 83.311 73.227 ;
      RECT 83.303 65.764 83.357 73.181 ;
      RECT 83.349 65.718 83.403 73.135 ;
      RECT 83.395 65.672 83.449 73.089 ;
      RECT 83.441 65.626 83.495 73.043 ;
      RECT 83.487 65.58 83.541 72.997 ;
      RECT 83.533 65.534 83.587 72.951 ;
      RECT 83.579 65.488 83.633 72.905 ;
      RECT 83.625 65.442 83.679 72.859 ;
      RECT 83.671 65.396 83.725 72.813 ;
      RECT 83.717 65.35 83.771 72.767 ;
      RECT 83.763 65.304 83.817 72.721 ;
      RECT 83.809 65.258 83.863 72.675 ;
      RECT 83.855 65.212 83.909 72.629 ;
      RECT 83.901 65.166 83.955 72.583 ;
      RECT 83.947 65.12 84.001 72.537 ;
      RECT 83.993 65.074 84.047 72.491 ;
      RECT 84.039 65.028 84.093 72.445 ;
      RECT 84.085 64.982 84.139 72.399 ;
      RECT 84.131 64.936 84.185 72.353 ;
      RECT 84.177 64.89 84.231 72.307 ;
      RECT 84.223 64.844 84.277 72.261 ;
      RECT 84.269 64.798 84.323 72.215 ;
      RECT 84.315 64.752 84.369 72.169 ;
      RECT 84.361 64.706 84.415 72.123 ;
      RECT 84.407 64.66 84.461 72.077 ;
      RECT 84.453 64.614 84.507 72.031 ;
      RECT 84.499 64.568 84.553 71.985 ;
      RECT 84.545 64.522 84.599 71.939 ;
      RECT 84.591 64.476 84.645 71.893 ;
      RECT 84.637 64.43 84.691 71.847 ;
      RECT 84.683 64.384 84.737 71.801 ;
      RECT 84.729 64.338 84.783 71.755 ;
      RECT 84.775 64.292 84.829 71.709 ;
      RECT 84.821 64.246 84.875 71.663 ;
      RECT 84.867 64.2 84.921 71.617 ;
      RECT 84.913 64.154 84.967 71.571 ;
      RECT 84.959 64.108 85.013 71.525 ;
      RECT 85.005 64.062 85.059 71.479 ;
      RECT 85.051 64.016 85.105 71.433 ;
      RECT 85.097 63.97 85.151 71.387 ;
      RECT 85.143 63.924 85.197 71.341 ;
      RECT 85.189 63.878 85.243 71.295 ;
      RECT 85.235 63.832 85.289 71.249 ;
      RECT 85.281 63.786 85.335 71.203 ;
      RECT 85.327 63.74 85.381 71.157 ;
      RECT 85.373 63.696 85.427 71.111 ;
      RECT 85.415 63.675 85.473 71.065 ;
      RECT 82.857 66.21 82.943 73.595 ;
      RECT 85.415 63.675 85.519 71.019 ;
      RECT 85.415 63.675 85.565 70.973 ;
      RECT 85.415 63.675 85.611 70.927 ;
      RECT 85.415 63.675 85.657 70.881 ;
      RECT 85.415 63.675 85.703 70.835 ;
      RECT 85.415 63.675 85.749 70.789 ;
      RECT 85.415 63.675 85.795 70.743 ;
      RECT 85.415 63.675 85.841 70.697 ;
      RECT 85.415 63.675 85.887 70.651 ;
      RECT 85.415 63.675 85.933 70.605 ;
      RECT 85.415 63.675 85.979 70.559 ;
      RECT 85.415 63.675 86.025 70.513 ;
      RECT 85.415 63.675 86.071 70.467 ;
      RECT 85.415 63.675 86.117 70.421 ;
      RECT 85.415 63.675 86.163 70.375 ;
      RECT 85.415 63.675 86.209 70.329 ;
      RECT 85.415 63.675 86.255 70.283 ;
      RECT 85.415 63.675 86.301 70.237 ;
      RECT 85.415 63.675 86.347 70.191 ;
      RECT 85.415 63.675 86.393 70.145 ;
      RECT 85.415 63.675 86.439 70.099 ;
      RECT 85.415 63.675 86.485 70.053 ;
      RECT 85.415 63.675 86.531 70.007 ;
      RECT 85.415 63.675 86.577 69.961 ;
      RECT 85.415 63.675 86.623 69.915 ;
      RECT 85.415 63.675 86.669 69.869 ;
      RECT 85.415 63.675 86.715 69.823 ;
      RECT 85.415 63.675 86.761 69.777 ;
      RECT 85.415 63.675 86.807 69.731 ;
      RECT 85.415 63.675 86.853 69.685 ;
      RECT 85.415 63.675 86.899 69.639 ;
      RECT 85.415 63.675 86.945 69.593 ;
      RECT 85.415 63.675 86.991 69.547 ;
      RECT 85.415 63.675 87.037 69.501 ;
      RECT 85.415 63.675 87.083 69.455 ;
      RECT 85.415 63.675 87.129 69.409 ;
      RECT 85.415 63.675 87.175 69.363 ;
      RECT 85.415 63.675 87.221 69.317 ;
      RECT 85.415 63.675 87.267 69.271 ;
      RECT 85.415 63.675 87.313 69.225 ;
      RECT 85.415 63.675 87.359 69.179 ;
      RECT 85.415 63.675 87.405 69.133 ;
      RECT 85.415 63.675 87.451 69.087 ;
      RECT 85.415 63.675 87.497 69.041 ;
      RECT 85.415 63.675 87.543 68.995 ;
      RECT 85.415 63.675 87.589 68.949 ;
      RECT 85.415 63.675 87.635 68.903 ;
      RECT 85.415 63.675 87.681 68.857 ;
      RECT 85.415 63.675 87.727 68.811 ;
      RECT 85.415 63.675 87.773 68.765 ;
      RECT 85.415 63.675 87.819 68.719 ;
      RECT 85.415 63.675 87.865 68.673 ;
      RECT 85.415 63.675 87.911 68.627 ;
      RECT 85.415 63.675 87.957 68.581 ;
      RECT 85.415 63.675 88.003 68.535 ;
      RECT 85.415 63.675 88.049 68.489 ;
      RECT 85.415 63.675 88.095 68.443 ;
      RECT 85.415 63.675 88.141 68.397 ;
      RECT 80.741 68.326 88.187 68.351 ;
      RECT 85.415 63.675 88.19 68.326 ;
      RECT 85.415 63.675 110 68.325 ;
      RECT 77.175 92.037 78.325 110 ;
      RECT 77.175 92.037 78.371 92.272 ;
      RECT 77.175 92.037 78.417 92.226 ;
      RECT 77.175 92.037 78.463 92.18 ;
      RECT 77.175 92.037 78.509 92.134 ;
      RECT 77.175 92.037 78.555 92.088 ;
      RECT 77.221 91.991 78.601 92.042 ;
      RECT 77.267 91.945 78.647 91.996 ;
      RECT 77.313 91.899 78.693 91.95 ;
      RECT 77.359 91.853 78.739 91.904 ;
      RECT 77.405 91.807 78.785 91.858 ;
      RECT 77.451 91.761 78.831 91.812 ;
      RECT 77.497 91.715 78.877 91.766 ;
      RECT 77.543 91.669 78.923 91.72 ;
      RECT 77.589 91.623 78.969 91.674 ;
      RECT 77.635 91.577 79.015 91.628 ;
      RECT 77.681 91.531 79.061 91.582 ;
      RECT 77.727 91.485 79.107 91.536 ;
      RECT 77.773 91.439 79.153 91.49 ;
      RECT 77.819 91.393 79.199 91.444 ;
      RECT 77.865 91.347 79.245 91.398 ;
      RECT 77.911 91.301 79.291 91.352 ;
      RECT 77.957 91.255 79.337 91.306 ;
      RECT 78.003 91.209 79.383 91.26 ;
      RECT 78.049 91.163 79.429 91.214 ;
      RECT 78.095 91.117 79.475 91.168 ;
      RECT 78.141 91.071 79.521 91.122 ;
      RECT 78.187 91.025 79.567 91.076 ;
      RECT 78.233 90.979 79.613 91.03 ;
      RECT 78.279 90.933 79.659 90.984 ;
      RECT 78.325 90.887 79.705 90.938 ;
      RECT 78.371 90.841 79.751 90.892 ;
      RECT 78.417 90.795 79.797 90.846 ;
      RECT 78.463 90.749 79.843 90.8 ;
      RECT 78.509 90.703 79.889 90.754 ;
      RECT 78.555 90.657 79.935 90.708 ;
      RECT 78.601 90.611 79.981 90.662 ;
      RECT 78.647 90.565 80.027 90.616 ;
      RECT 78.693 90.519 80.073 90.57 ;
      RECT 78.739 90.473 80.119 90.524 ;
      RECT 78.785 90.427 80.165 90.478 ;
      RECT 78.831 90.381 80.211 90.432 ;
      RECT 78.877 90.335 80.257 90.386 ;
      RECT 78.923 90.289 80.303 90.34 ;
      RECT 78.969 90.243 80.349 90.294 ;
      RECT 79.015 90.197 80.395 90.248 ;
      RECT 79.061 90.151 80.441 90.202 ;
      RECT 79.107 90.105 80.487 90.156 ;
      RECT 79.153 90.059 80.533 90.11 ;
      RECT 79.199 90.013 80.579 90.064 ;
      RECT 79.245 89.967 80.625 90.018 ;
      RECT 79.291 89.921 80.671 89.972 ;
      RECT 79.337 89.875 80.717 89.926 ;
      RECT 79.383 89.829 80.763 89.88 ;
      RECT 79.429 89.783 80.809 89.834 ;
      RECT 79.475 89.737 80.855 89.788 ;
      RECT 79.521 89.691 80.901 89.742 ;
      RECT 79.567 89.645 80.947 89.696 ;
      RECT 79.613 89.599 80.993 89.65 ;
      RECT 79.659 89.553 81.039 89.604 ;
      RECT 79.705 89.507 81.085 89.558 ;
      RECT 79.751 89.461 81.131 89.512 ;
      RECT 79.797 89.415 81.177 89.466 ;
      RECT 79.843 89.369 81.223 89.42 ;
      RECT 79.889 89.323 81.269 89.374 ;
      RECT 79.935 89.277 81.315 89.328 ;
      RECT 79.981 89.231 81.361 89.282 ;
      RECT 80.027 89.185 81.407 89.236 ;
      RECT 80.073 89.139 81.453 89.19 ;
      RECT 80.119 89.093 81.499 89.144 ;
      RECT 80.165 89.047 81.545 89.098 ;
      RECT 80.211 89.001 81.591 89.052 ;
      RECT 80.257 88.955 81.637 89.006 ;
      RECT 80.303 88.909 81.683 88.96 ;
      RECT 80.349 88.863 81.729 88.914 ;
      RECT 80.395 88.817 81.775 88.868 ;
      RECT 80.441 88.771 81.821 88.822 ;
      RECT 80.487 88.725 81.867 88.776 ;
      RECT 80.533 88.679 81.913 88.73 ;
      RECT 80.579 88.633 81.959 88.684 ;
      RECT 80.625 88.587 82.005 88.638 ;
      RECT 80.671 88.541 82.051 88.592 ;
      RECT 80.717 88.495 82.097 88.546 ;
      RECT 80.763 88.449 82.143 88.5 ;
      RECT 80.809 88.403 82.189 88.454 ;
      RECT 80.855 88.357 82.235 88.408 ;
      RECT 80.901 88.311 82.281 88.362 ;
      RECT 80.947 88.265 82.327 88.316 ;
      RECT 80.993 88.219 82.373 88.27 ;
      RECT 81.039 88.173 82.419 88.224 ;
      RECT 81.085 88.127 82.465 88.178 ;
      RECT 81.131 88.081 82.511 88.132 ;
      RECT 81.177 88.035 82.557 88.086 ;
      RECT 81.223 87.989 82.603 88.04 ;
      RECT 81.269 87.943 82.649 87.994 ;
      RECT 81.315 87.897 82.695 87.948 ;
      RECT 81.361 87.851 82.741 87.902 ;
      RECT 81.407 87.805 82.787 87.856 ;
      RECT 81.453 87.759 82.833 87.81 ;
      RECT 81.499 87.713 82.879 87.764 ;
      RECT 81.545 87.667 82.925 87.718 ;
      RECT 81.591 87.621 82.971 87.672 ;
      RECT 81.637 87.575 83.017 87.626 ;
      RECT 81.683 87.529 83.063 87.58 ;
      RECT 81.729 87.483 83.109 87.534 ;
      RECT 81.775 87.437 83.155 87.488 ;
      RECT 81.821 87.391 83.201 87.442 ;
      RECT 81.867 87.345 83.247 87.396 ;
      RECT 81.913 87.299 83.293 87.35 ;
      RECT 81.959 87.253 83.339 87.304 ;
      RECT 82.005 87.207 83.385 87.258 ;
      RECT 82.051 87.161 83.431 87.212 ;
      RECT 82.097 87.115 83.477 87.166 ;
      RECT 82.143 87.069 83.523 87.12 ;
      RECT 82.189 87.023 83.569 87.074 ;
      RECT 82.235 86.977 83.615 87.028 ;
      RECT 82.281 86.931 83.661 86.982 ;
      RECT 82.327 86.885 83.707 86.936 ;
      RECT 82.373 86.839 83.753 86.89 ;
      RECT 82.419 86.793 83.799 86.844 ;
      RECT 82.465 86.747 83.845 86.798 ;
      RECT 82.511 86.701 83.891 86.752 ;
      RECT 82.557 86.655 83.937 86.706 ;
      RECT 82.603 86.609 83.983 86.66 ;
      RECT 82.649 86.563 84.029 86.614 ;
      RECT 82.695 86.517 84.075 86.568 ;
      RECT 82.741 86.471 84.121 86.522 ;
      RECT 82.787 86.425 84.167 86.476 ;
      RECT 82.833 86.379 84.213 86.43 ;
      RECT 82.879 86.333 84.259 86.384 ;
      RECT 82.925 86.287 84.305 86.338 ;
      RECT 82.971 86.241 84.351 86.292 ;
      RECT 83.017 86.195 84.397 86.246 ;
      RECT 83.063 86.149 84.443 86.2 ;
      RECT 83.109 86.103 84.489 86.154 ;
      RECT 83.155 86.057 84.535 86.108 ;
      RECT 83.201 86.011 84.581 86.062 ;
      RECT 83.247 85.965 84.627 86.016 ;
      RECT 83.293 85.919 84.673 85.97 ;
      RECT 83.339 85.873 84.719 85.924 ;
      RECT 83.385 85.827 84.765 85.878 ;
      RECT 83.431 85.781 84.811 85.832 ;
      RECT 83.477 85.735 84.857 85.786 ;
      RECT 83.523 85.689 84.903 85.74 ;
      RECT 83.569 85.643 84.949 85.694 ;
      RECT 83.615 85.597 84.995 85.648 ;
      RECT 83.661 85.551 85.041 85.602 ;
      RECT 83.707 85.505 85.087 85.556 ;
      RECT 83.753 85.459 85.133 85.51 ;
      RECT 83.799 85.413 85.179 85.464 ;
      RECT 83.845 85.367 85.225 85.418 ;
      RECT 83.891 85.321 85.271 85.372 ;
      RECT 83.937 85.275 85.317 85.326 ;
      RECT 83.983 85.229 85.363 85.28 ;
      RECT 84.029 85.183 85.409 85.234 ;
      RECT 84.075 85.137 85.455 85.188 ;
      RECT 84.121 85.091 85.501 85.142 ;
      RECT 84.167 85.045 85.547 85.096 ;
      RECT 84.213 84.999 85.593 85.05 ;
      RECT 84.259 84.953 85.639 85.004 ;
      RECT 84.305 84.907 85.685 84.958 ;
      RECT 84.351 84.861 85.731 84.912 ;
      RECT 84.397 84.815 85.777 84.866 ;
      RECT 84.443 84.769 85.823 84.82 ;
      RECT 84.489 84.723 85.869 84.774 ;
      RECT 84.535 84.677 85.915 84.728 ;
      RECT 84.581 84.631 85.961 84.682 ;
      RECT 84.627 84.585 86.007 84.636 ;
      RECT 84.673 84.539 86.053 84.59 ;
      RECT 84.719 84.493 86.099 84.544 ;
      RECT 84.765 84.447 86.145 84.498 ;
      RECT 84.811 84.401 86.191 84.452 ;
      RECT 84.857 84.355 86.237 84.406 ;
      RECT 84.903 84.309 86.283 84.36 ;
      RECT 84.949 84.263 86.329 84.314 ;
      RECT 84.995 84.217 86.375 84.268 ;
      RECT 85.041 84.171 86.421 84.222 ;
      RECT 85.087 84.125 86.467 84.176 ;
      RECT 85.133 84.079 86.513 84.13 ;
      RECT 85.179 84.033 86.559 84.084 ;
      RECT 85.225 83.987 86.605 84.038 ;
      RECT 85.271 83.941 86.651 83.992 ;
      RECT 85.317 83.895 86.697 83.946 ;
      RECT 85.363 83.849 86.743 83.9 ;
      RECT 85.409 83.803 86.789 83.854 ;
      RECT 85.455 83.757 86.835 83.808 ;
      RECT 85.501 83.711 86.881 83.762 ;
      RECT 85.547 83.665 86.927 83.716 ;
      RECT 85.593 83.619 86.973 83.67 ;
      RECT 85.639 83.573 87.019 83.624 ;
      RECT 85.685 83.527 87.065 83.578 ;
      RECT 85.731 83.481 87.111 83.532 ;
      RECT 85.777 83.435 87.157 83.486 ;
      RECT 85.823 83.389 87.203 83.44 ;
      RECT 85.869 83.343 87.249 83.394 ;
      RECT 85.915 83.297 87.295 83.348 ;
      RECT 85.961 83.251 87.341 83.302 ;
      RECT 86.007 83.205 87.387 83.256 ;
      RECT 86.053 83.159 87.433 83.21 ;
      RECT 86.099 83.113 87.479 83.164 ;
      RECT 86.145 83.067 87.525 83.118 ;
      RECT 86.191 83.021 87.571 83.072 ;
      RECT 86.237 82.975 87.617 83.026 ;
      RECT 86.283 82.929 87.663 82.98 ;
      RECT 86.329 82.883 87.709 82.934 ;
      RECT 86.375 82.837 87.755 82.888 ;
      RECT 86.421 82.791 87.801 82.842 ;
      RECT 86.467 82.745 87.847 82.796 ;
      RECT 86.513 82.699 87.893 82.75 ;
      RECT 86.559 82.653 87.939 82.704 ;
      RECT 86.605 82.607 87.985 82.658 ;
      RECT 86.651 82.561 88.031 82.612 ;
      RECT 86.697 82.515 88.077 82.566 ;
      RECT 86.743 82.469 88.123 82.52 ;
      RECT 86.789 82.423 88.169 82.474 ;
      RECT 86.835 82.377 88.215 82.428 ;
      RECT 86.881 82.331 88.261 82.382 ;
      RECT 86.927 82.285 88.307 82.336 ;
      RECT 86.973 82.239 88.353 82.29 ;
      RECT 87.019 82.193 88.399 82.244 ;
      RECT 87.065 82.147 88.445 82.198 ;
      RECT 87.111 82.101 88.491 82.152 ;
      RECT 87.157 82.055 88.537 82.106 ;
      RECT 87.203 82.009 88.583 82.06 ;
      RECT 88.537 80.697 88.583 82.06 ;
      RECT 87.249 81.963 88.629 82.014 ;
      RECT 87.295 81.917 88.675 81.968 ;
      RECT 87.341 81.871 88.721 81.922 ;
      RECT 87.387 81.825 88.767 81.876 ;
      RECT 87.433 81.779 88.813 81.83 ;
      RECT 87.479 81.733 88.859 81.784 ;
      RECT 87.525 81.687 88.905 81.738 ;
      RECT 87.571 81.641 88.951 81.692 ;
      RECT 87.617 81.595 88.997 81.646 ;
      RECT 87.663 81.549 89.043 81.6 ;
      RECT 87.709 81.503 89.089 81.554 ;
      RECT 87.755 81.457 89.135 81.508 ;
      RECT 87.801 81.411 89.181 81.462 ;
      RECT 87.847 81.365 89.227 81.416 ;
      RECT 87.893 81.319 89.273 81.37 ;
      RECT 87.939 81.273 89.319 81.324 ;
      RECT 87.939 81.273 89.325 81.298 ;
      RECT 87.985 81.227 89.371 81.272 ;
      RECT 88.031 81.181 89.417 81.226 ;
      RECT 88.077 81.135 89.463 81.18 ;
      RECT 88.123 81.089 89.509 81.134 ;
      RECT 88.169 81.043 89.555 81.088 ;
      RECT 88.215 80.997 89.601 81.042 ;
      RECT 88.261 80.951 89.647 80.996 ;
      RECT 88.307 80.905 89.693 80.95 ;
      RECT 88.353 80.859 89.739 80.904 ;
      RECT 88.399 80.813 89.785 80.858 ;
      RECT 88.445 80.767 89.831 80.812 ;
      RECT 88.491 80.721 89.877 80.766 ;
      RECT 88.54 80.672 89.923 80.72 ;
      RECT 89.874 79.338 89.923 80.72 ;
      RECT 88.586 80.626 89.969 80.674 ;
      RECT 89.92 79.292 89.969 80.674 ;
      RECT 88.632 80.58 90.015 80.628 ;
      RECT 89.966 79.246 90.015 80.628 ;
      RECT 88.678 80.534 90.061 80.582 ;
      RECT 90.012 79.2 90.061 80.582 ;
      RECT 88.724 80.488 90.107 80.536 ;
      RECT 90.058 79.154 90.107 80.536 ;
      RECT 88.77 80.442 90.153 80.49 ;
      RECT 90.104 79.108 90.153 80.49 ;
      RECT 88.816 80.396 90.199 80.444 ;
      RECT 90.15 79.062 90.199 80.444 ;
      RECT 88.862 80.35 90.245 80.398 ;
      RECT 90.196 79.016 90.245 80.398 ;
      RECT 88.908 80.304 90.291 80.352 ;
      RECT 90.242 78.97 90.291 80.352 ;
      RECT 88.954 80.258 90.337 80.306 ;
      RECT 90.288 78.924 90.337 80.306 ;
      RECT 89 80.212 90.383 80.26 ;
      RECT 90.334 78.878 90.383 80.26 ;
      RECT 89.046 80.166 90.429 80.214 ;
      RECT 90.38 78.832 90.429 80.214 ;
      RECT 89.092 80.12 90.475 80.168 ;
      RECT 90.426 78.786 90.475 80.168 ;
      RECT 89.138 80.074 90.521 80.122 ;
      RECT 90.472 78.74 90.521 80.122 ;
      RECT 89.184 80.028 90.567 80.076 ;
      RECT 90.518 78.694 90.567 80.076 ;
      RECT 89.23 79.982 90.613 80.03 ;
      RECT 90.564 78.648 90.613 80.03 ;
      RECT 89.276 79.936 90.659 79.984 ;
      RECT 90.61 78.602 90.659 79.984 ;
      RECT 89.322 79.89 90.705 79.938 ;
      RECT 90.656 78.556 90.705 79.938 ;
      RECT 89.368 79.844 90.751 79.892 ;
      RECT 90.702 78.51 90.751 79.892 ;
      RECT 89.414 79.798 90.797 79.846 ;
      RECT 90.748 78.464 90.797 79.846 ;
      RECT 89.46 79.752 90.843 79.8 ;
      RECT 90.794 78.418 90.843 79.8 ;
      RECT 89.506 79.706 90.889 79.754 ;
      RECT 90.84 78.372 90.889 79.754 ;
      RECT 89.552 79.66 90.935 79.708 ;
      RECT 90.886 78.326 90.935 79.708 ;
      RECT 89.598 79.614 90.981 79.662 ;
      RECT 90.932 78.28 90.981 79.662 ;
      RECT 89.644 79.568 91.027 79.616 ;
      RECT 90.978 78.234 91.027 79.616 ;
      RECT 89.69 79.522 91.073 79.57 ;
      RECT 91.024 78.188 91.073 79.57 ;
      RECT 89.736 79.476 91.119 79.524 ;
      RECT 91.07 78.142 91.119 79.524 ;
      RECT 89.782 79.43 91.165 79.478 ;
      RECT 91.116 78.096 91.165 79.478 ;
      RECT 89.828 79.384 91.211 79.432 ;
      RECT 91.162 78.05 91.211 79.432 ;
      RECT 91.208 78.004 91.257 79.386 ;
      RECT 91.254 77.958 91.303 79.34 ;
      RECT 91.3 77.912 91.349 79.294 ;
      RECT 91.346 77.866 91.395 79.248 ;
      RECT 91.392 77.82 91.441 79.202 ;
      RECT 91.438 77.774 91.487 79.156 ;
      RECT 91.484 77.728 91.533 79.11 ;
      RECT 91.53 77.682 91.579 79.064 ;
      RECT 91.576 77.636 91.625 79.018 ;
      RECT 91.622 77.59 91.671 78.972 ;
      RECT 91.668 77.544 91.717 78.926 ;
      RECT 91.714 77.498 91.763 78.88 ;
      RECT 91.76 77.452 91.809 78.834 ;
      RECT 91.806 77.406 91.855 78.788 ;
      RECT 91.852 77.36 91.901 78.742 ;
      RECT 91.898 77.314 91.947 78.696 ;
      RECT 91.944 77.268 91.993 78.65 ;
      RECT 91.99 77.222 92.039 78.604 ;
      RECT 92.036 77.187 92.085 78.558 ;
      RECT 92.06 77.175 92.131 78.512 ;
      RECT 92.06 77.175 92.177 78.466 ;
      RECT 92.06 77.175 92.223 78.42 ;
      RECT 92.06 77.175 92.269 78.374 ;
      RECT 90.886 78.326 92.295 78.338 ;
      RECT 92.06 77.175 110 78.325 ;
      RECT 89.675 97.182 90.825 110 ;
      RECT 89.675 97.182 90.871 99.352 ;
      RECT 89.675 97.182 90.917 99.306 ;
      RECT 89.675 97.182 90.963 99.26 ;
      RECT 89.675 97.182 91.009 99.214 ;
      RECT 89.675 97.182 91.055 99.168 ;
      RECT 89.675 97.182 91.101 99.122 ;
      RECT 89.675 97.182 91.147 99.076 ;
      RECT 89.675 97.182 91.193 99.03 ;
      RECT 89.675 97.182 91.239 98.984 ;
      RECT 89.675 97.182 91.285 98.938 ;
      RECT 89.675 97.182 91.331 98.892 ;
      RECT 89.675 97.182 91.377 98.846 ;
      RECT 89.675 97.182 91.423 98.8 ;
      RECT 89.675 97.182 91.469 98.754 ;
      RECT 89.675 97.182 91.515 98.708 ;
      RECT 89.675 97.182 91.561 98.662 ;
      RECT 89.675 97.182 91.607 98.616 ;
      RECT 89.675 97.182 91.653 98.57 ;
      RECT 89.675 97.182 91.699 98.524 ;
      RECT 89.675 97.182 91.745 98.478 ;
      RECT 89.675 97.182 91.791 98.432 ;
      RECT 89.675 97.182 91.837 98.386 ;
      RECT 89.675 97.182 91.883 98.34 ;
      RECT 89.675 97.182 91.929 98.294 ;
      RECT 89.675 97.182 91.975 98.248 ;
      RECT 89.675 97.182 92.021 98.202 ;
      RECT 89.675 97.182 92.067 98.156 ;
      RECT 89.675 97.182 92.113 98.11 ;
      RECT 89.675 97.182 92.159 98.064 ;
      RECT 89.675 97.182 92.205 98.018 ;
      RECT 89.675 97.182 92.251 97.972 ;
      RECT 89.675 97.182 92.297 97.926 ;
      RECT 89.675 97.182 92.343 97.88 ;
      RECT 89.675 97.182 92.389 97.834 ;
      RECT 89.675 97.182 92.435 97.788 ;
      RECT 89.675 97.182 92.481 97.742 ;
      RECT 89.675 97.182 92.527 97.696 ;
      RECT 89.675 97.182 92.573 97.65 ;
      RECT 89.675 97.182 92.619 97.604 ;
      RECT 89.675 97.182 92.665 97.558 ;
      RECT 89.675 97.182 92.711 97.512 ;
      RECT 89.675 97.182 92.757 97.466 ;
      RECT 89.675 97.182 92.803 97.42 ;
      RECT 89.675 97.182 92.849 97.374 ;
      RECT 89.675 97.182 92.895 97.328 ;
      RECT 89.675 97.182 92.941 97.282 ;
      RECT 89.721 97.136 93.033 97.19 ;
      RECT 92.967 93.89 93.033 97.19 ;
      RECT 89.767 97.09 93.079 97.144 ;
      RECT 93.013 93.844 93.079 97.144 ;
      RECT 89.813 97.044 93.125 97.098 ;
      RECT 93.059 93.798 93.125 97.098 ;
      RECT 89.859 96.998 93.171 97.052 ;
      RECT 93.105 93.752 93.171 97.052 ;
      RECT 89.905 96.952 93.217 97.006 ;
      RECT 93.151 93.706 93.217 97.006 ;
      RECT 89.951 96.906 93.263 96.96 ;
      RECT 93.197 93.66 93.263 96.96 ;
      RECT 89.997 96.86 93.309 96.914 ;
      RECT 93.243 93.614 93.309 96.914 ;
      RECT 90.043 96.814 93.355 96.868 ;
      RECT 93.289 93.568 93.355 96.868 ;
      RECT 90.089 96.768 93.401 96.822 ;
      RECT 93.335 93.522 93.401 96.822 ;
      RECT 90.135 96.722 93.447 96.776 ;
      RECT 93.381 93.476 93.447 96.776 ;
      RECT 90.181 96.676 93.493 96.73 ;
      RECT 93.427 93.43 93.493 96.73 ;
      RECT 90.227 96.63 93.539 96.684 ;
      RECT 93.473 93.384 93.539 96.684 ;
      RECT 90.273 96.584 93.585 96.638 ;
      RECT 93.519 93.338 93.585 96.638 ;
      RECT 90.319 96.538 93.631 96.592 ;
      RECT 93.565 93.292 93.631 96.592 ;
      RECT 90.365 96.492 93.677 96.546 ;
      RECT 93.611 93.246 93.677 96.546 ;
      RECT 90.411 96.446 93.723 96.5 ;
      RECT 93.657 93.2 93.723 96.5 ;
      RECT 90.457 96.4 93.769 96.454 ;
      RECT 93.703 93.154 93.769 96.454 ;
      RECT 90.503 96.354 93.815 96.408 ;
      RECT 93.749 93.108 93.815 96.408 ;
      RECT 90.549 96.308 93.861 96.362 ;
      RECT 93.795 93.062 93.861 96.362 ;
      RECT 90.595 96.262 93.907 96.316 ;
      RECT 93.841 93.016 93.907 96.316 ;
      RECT 90.641 96.216 93.953 96.27 ;
      RECT 93.887 92.97 93.953 96.27 ;
      RECT 90.687 96.17 93.999 96.224 ;
      RECT 93.933 92.924 93.999 96.224 ;
      RECT 90.733 96.124 94.045 96.178 ;
      RECT 93.979 92.878 94.045 96.178 ;
      RECT 90.779 96.078 94.091 96.132 ;
      RECT 94.025 92.832 94.091 96.132 ;
      RECT 90.825 96.032 94.137 96.086 ;
      RECT 94.071 92.786 94.137 96.086 ;
      RECT 90.871 95.986 94.183 96.04 ;
      RECT 94.117 92.74 94.183 96.04 ;
      RECT 90.917 95.94 94.229 95.994 ;
      RECT 94.163 92.694 94.229 95.994 ;
      RECT 90.963 95.894 94.275 95.948 ;
      RECT 94.209 92.648 94.275 95.948 ;
      RECT 91.009 95.848 94.321 95.902 ;
      RECT 94.255 92.602 94.321 95.902 ;
      RECT 91.055 95.802 94.367 95.856 ;
      RECT 94.301 92.556 94.367 95.856 ;
      RECT 91.101 95.756 94.413 95.81 ;
      RECT 94.347 92.51 94.413 95.81 ;
      RECT 91.147 95.71 94.459 95.764 ;
      RECT 94.393 92.464 94.459 95.764 ;
      RECT 91.193 95.664 94.505 95.718 ;
      RECT 94.439 92.418 94.505 95.718 ;
      RECT 91.239 95.618 94.551 95.672 ;
      RECT 94.485 92.372 94.551 95.672 ;
      RECT 91.285 95.572 94.597 95.626 ;
      RECT 94.531 92.326 94.597 95.626 ;
      RECT 91.331 95.526 94.643 95.58 ;
      RECT 94.577 92.28 94.643 95.58 ;
      RECT 91.377 95.48 94.689 95.534 ;
      RECT 94.623 92.234 94.689 95.534 ;
      RECT 91.423 95.434 94.735 95.488 ;
      RECT 94.669 92.188 94.735 95.488 ;
      RECT 91.469 95.388 94.781 95.442 ;
      RECT 94.715 92.142 94.781 95.442 ;
      RECT 91.515 95.342 94.827 95.396 ;
      RECT 94.761 92.096 94.827 95.396 ;
      RECT 91.561 95.296 94.873 95.35 ;
      RECT 94.807 92.05 94.873 95.35 ;
      RECT 91.607 95.25 94.919 95.304 ;
      RECT 94.853 92.004 94.919 95.304 ;
      RECT 91.653 95.204 94.965 95.258 ;
      RECT 94.899 91.958 94.965 95.258 ;
      RECT 91.699 95.158 95.011 95.212 ;
      RECT 94.945 91.912 95.011 95.212 ;
      RECT 91.745 95.112 95.057 95.166 ;
      RECT 94.991 91.866 95.057 95.166 ;
      RECT 91.791 95.066 95.103 95.12 ;
      RECT 95.037 91.82 95.103 95.12 ;
      RECT 91.837 95.02 95.149 95.074 ;
      RECT 95.083 91.774 95.149 95.074 ;
      RECT 91.883 94.974 95.195 95.028 ;
      RECT 95.129 91.728 95.195 95.028 ;
      RECT 91.929 94.928 95.241 94.982 ;
      RECT 95.175 91.682 95.241 94.982 ;
      RECT 91.975 94.882 95.287 94.936 ;
      RECT 95.221 91.636 95.287 94.936 ;
      RECT 92.021 94.836 95.333 94.89 ;
      RECT 95.267 91.59 95.333 94.89 ;
      RECT 92.067 94.79 95.379 94.844 ;
      RECT 95.313 91.544 95.379 94.844 ;
      RECT 92.113 94.744 95.425 94.798 ;
      RECT 95.359 91.498 95.425 94.798 ;
      RECT 92.159 94.698 95.471 94.752 ;
      RECT 95.405 91.452 95.471 94.752 ;
      RECT 92.205 94.652 95.517 94.706 ;
      RECT 95.451 91.406 95.517 94.706 ;
      RECT 92.251 94.606 95.563 94.66 ;
      RECT 95.497 91.36 95.563 94.66 ;
      RECT 92.297 94.56 95.609 94.614 ;
      RECT 95.543 91.314 95.609 94.614 ;
      RECT 92.343 94.514 95.655 94.568 ;
      RECT 95.589 91.268 95.655 94.568 ;
      RECT 92.389 94.468 95.701 94.522 ;
      RECT 95.635 91.222 95.701 94.522 ;
      RECT 92.435 94.422 95.747 94.476 ;
      RECT 95.681 91.176 95.747 94.476 ;
      RECT 92.481 94.376 95.793 94.43 ;
      RECT 95.727 91.13 95.793 94.43 ;
      RECT 92.527 94.33 95.839 94.384 ;
      RECT 95.773 91.084 95.839 94.384 ;
      RECT 92.573 94.284 95.885 94.338 ;
      RECT 95.819 91.038 95.885 94.338 ;
      RECT 92.619 94.248 95.931 94.292 ;
      RECT 95.865 90.992 95.931 94.292 ;
      RECT 92.645 94.212 95.931 94.292 ;
      RECT 92.921 93.936 92.987 97.236 ;
      RECT 92.691 94.166 95.977 94.246 ;
      RECT 95.911 90.946 95.977 94.246 ;
      RECT 92.737 94.12 96.023 94.2 ;
      RECT 95.957 90.9 96.023 94.2 ;
      RECT 92.783 94.074 96.069 94.154 ;
      RECT 96.003 90.854 96.069 94.154 ;
      RECT 92.829 94.028 96.115 94.108 ;
      RECT 96.049 90.808 96.115 94.108 ;
      RECT 92.875 93.982 96.161 94.062 ;
      RECT 96.095 90.762 96.161 94.062 ;
      RECT 96.141 90.716 96.207 94.016 ;
      RECT 96.187 90.67 96.253 93.97 ;
      RECT 96.233 90.624 96.299 93.924 ;
      RECT 96.279 90.578 96.345 93.878 ;
      RECT 96.325 90.532 96.391 93.832 ;
      RECT 96.371 90.486 96.437 93.786 ;
      RECT 96.417 90.44 96.483 93.74 ;
      RECT 96.463 90.394 96.529 93.694 ;
      RECT 96.509 90.348 96.575 93.648 ;
      RECT 96.555 90.302 96.621 93.602 ;
      RECT 96.601 90.256 96.667 93.556 ;
      RECT 96.647 90.21 96.713 93.51 ;
      RECT 96.693 90.164 96.759 93.464 ;
      RECT 96.739 90.118 96.805 93.418 ;
      RECT 96.785 90.072 96.851 93.372 ;
      RECT 96.831 90.026 96.897 93.326 ;
      RECT 96.877 89.98 96.943 93.28 ;
      RECT 96.923 89.934 96.989 93.234 ;
      RECT 96.969 89.888 97.035 93.188 ;
      RECT 97.015 89.842 97.081 93.142 ;
      RECT 97.061 89.796 97.127 93.096 ;
      RECT 97.107 89.75 97.173 93.05 ;
      RECT 97.199 89.678 97.219 93.004 ;
      RECT 97.205 89.675 97.265 92.958 ;
      RECT 97.153 89.704 97.219 93.004 ;
      RECT 97.205 89.675 97.311 92.912 ;
      RECT 97.205 89.675 97.357 92.866 ;
      RECT 97.205 89.675 97.403 92.82 ;
      RECT 97.205 89.675 97.449 92.774 ;
      RECT 97.205 89.675 97.495 92.728 ;
      RECT 97.205 89.675 97.541 92.682 ;
      RECT 97.205 89.675 97.587 92.636 ;
      RECT 97.205 89.675 97.633 92.59 ;
      RECT 97.205 89.675 97.679 92.544 ;
      RECT 97.205 89.675 97.725 92.498 ;
      RECT 97.205 89.675 97.771 92.452 ;
      RECT 94.485 92.372 97.817 92.406 ;
      RECT 97.205 89.675 97.825 92.379 ;
      RECT 97.205 89.675 97.871 92.352 ;
      RECT 97.205 89.675 97.917 92.306 ;
      RECT 97.205 89.675 97.963 92.26 ;
      RECT 97.205 89.675 98.009 92.214 ;
      RECT 97.205 89.675 98.055 92.168 ;
      RECT 97.205 89.675 98.101 92.122 ;
      RECT 97.205 89.675 98.147 92.076 ;
      RECT 97.205 89.675 98.193 92.03 ;
      RECT 97.205 89.675 98.239 91.984 ;
      RECT 97.205 89.675 98.285 91.938 ;
      RECT 97.205 89.675 98.331 91.892 ;
      RECT 97.205 89.675 98.377 91.846 ;
      RECT 97.205 89.675 98.423 91.8 ;
      RECT 97.205 89.675 98.469 91.754 ;
      RECT 97.205 89.675 98.515 91.708 ;
      RECT 97.205 89.675 98.561 91.662 ;
      RECT 97.205 89.675 98.607 91.616 ;
      RECT 97.205 89.675 98.653 91.57 ;
      RECT 97.205 89.675 98.699 91.524 ;
      RECT 97.205 89.675 98.745 91.478 ;
      RECT 97.205 89.675 98.791 91.432 ;
      RECT 97.205 89.675 98.837 91.386 ;
      RECT 97.205 89.675 98.883 91.34 ;
      RECT 97.205 89.675 98.929 91.294 ;
      RECT 97.205 89.675 98.975 91.248 ;
      RECT 97.205 89.675 99.021 91.202 ;
      RECT 97.205 89.675 99.067 91.156 ;
      RECT 97.205 89.675 99.113 91.11 ;
      RECT 97.205 89.675 99.159 91.064 ;
      RECT 97.205 89.675 99.205 91.018 ;
      RECT 97.205 89.675 99.251 90.972 ;
      RECT 97.205 89.675 99.297 90.926 ;
      RECT 97.205 89.675 99.343 90.88 ;
      RECT 96.049 90.808 99.375 90.841 ;
      RECT 97.205 89.675 110 90.825 ;
      RECT 98.175 102.602 99.325 110 ;
      RECT 98.175 102.602 99.371 103.642 ;
      RECT 98.175 102.602 99.417 103.596 ;
      RECT 98.175 102.602 99.463 103.55 ;
      RECT 98.175 102.602 99.509 103.504 ;
      RECT 98.175 102.602 99.555 103.458 ;
      RECT 98.175 102.602 99.601 103.412 ;
      RECT 98.175 102.602 99.647 103.366 ;
      RECT 98.175 102.602 99.693 103.32 ;
      RECT 98.175 102.602 99.739 103.274 ;
      RECT 98.175 102.602 99.785 103.228 ;
      RECT 98.175 102.602 99.831 103.182 ;
      RECT 98.175 102.602 99.877 103.136 ;
      RECT 98.175 102.602 99.923 103.09 ;
      RECT 98.175 102.602 99.969 103.044 ;
      RECT 98.175 102.602 100.015 102.998 ;
      RECT 98.175 102.602 100.061 102.952 ;
      RECT 98.175 102.602 100.107 102.906 ;
      RECT 98.175 102.602 100.153 102.86 ;
      RECT 98.175 102.602 100.199 102.814 ;
      RECT 98.175 102.602 100.245 102.768 ;
      RECT 98.175 102.602 100.291 102.722 ;
      RECT 98.175 102.602 100.337 102.676 ;
      RECT 98.221 102.556 100.383 102.63 ;
      RECT 100.323 100.454 100.383 102.63 ;
      RECT 98.267 102.51 100.429 102.584 ;
      RECT 100.369 100.408 100.429 102.584 ;
      RECT 98.313 102.464 100.475 102.538 ;
      RECT 100.415 100.362 100.475 102.538 ;
      RECT 98.359 102.418 100.521 102.492 ;
      RECT 100.461 100.316 100.521 102.492 ;
      RECT 98.405 102.372 100.567 102.446 ;
      RECT 100.507 100.27 100.567 102.446 ;
      RECT 98.451 102.326 100.613 102.4 ;
      RECT 100.553 100.224 100.613 102.4 ;
      RECT 98.497 102.28 100.659 102.354 ;
      RECT 100.599 100.178 100.659 102.354 ;
      RECT 98.543 102.234 100.705 102.308 ;
      RECT 100.645 100.132 100.705 102.308 ;
      RECT 98.589 102.188 100.751 102.262 ;
      RECT 100.691 100.086 100.751 102.262 ;
      RECT 98.635 102.142 100.797 102.216 ;
      RECT 100.737 100.04 100.797 102.216 ;
      RECT 98.681 102.096 100.843 102.17 ;
      RECT 100.783 99.994 100.843 102.17 ;
      RECT 98.727 102.05 100.889 102.124 ;
      RECT 100.829 99.948 100.889 102.124 ;
      RECT 98.773 102.004 100.935 102.078 ;
      RECT 100.875 99.902 100.935 102.078 ;
      RECT 98.819 101.958 100.981 102.032 ;
      RECT 100.921 99.856 100.981 102.032 ;
      RECT 98.865 101.912 101.027 101.986 ;
      RECT 100.967 99.81 101.027 101.986 ;
      RECT 98.911 101.866 101.073 101.94 ;
      RECT 101.013 99.764 101.073 101.94 ;
      RECT 98.957 101.82 101.119 101.894 ;
      RECT 101.059 99.718 101.119 101.894 ;
      RECT 99.003 101.774 101.165 101.848 ;
      RECT 101.105 99.672 101.165 101.848 ;
      RECT 99.049 101.728 101.211 101.802 ;
      RECT 101.151 99.626 101.211 101.802 ;
      RECT 99.095 101.682 101.257 101.756 ;
      RECT 101.197 99.58 101.257 101.756 ;
      RECT 99.141 101.636 101.303 101.71 ;
      RECT 101.243 99.534 101.303 101.71 ;
      RECT 99.187 101.59 101.349 101.664 ;
      RECT 101.289 99.488 101.349 101.664 ;
      RECT 99.233 101.544 101.395 101.618 ;
      RECT 101.335 99.442 101.395 101.618 ;
      RECT 99.279 101.498 101.441 101.572 ;
      RECT 101.381 99.396 101.441 101.572 ;
      RECT 99.325 101.452 101.487 101.526 ;
      RECT 101.427 99.35 101.487 101.526 ;
      RECT 99.371 101.406 101.533 101.48 ;
      RECT 101.473 99.304 101.533 101.48 ;
      RECT 99.417 101.36 101.579 101.434 ;
      RECT 101.519 99.258 101.579 101.434 ;
      RECT 99.463 101.314 101.625 101.388 ;
      RECT 101.565 99.212 101.625 101.388 ;
      RECT 99.509 101.268 101.671 101.342 ;
      RECT 101.611 99.166 101.671 101.342 ;
      RECT 99.555 101.222 101.717 101.296 ;
      RECT 101.657 99.12 101.717 101.296 ;
      RECT 99.601 101.176 101.763 101.25 ;
      RECT 101.703 99.074 101.763 101.25 ;
      RECT 99.647 101.13 101.809 101.204 ;
      RECT 101.749 99.028 101.809 101.204 ;
      RECT 99.693 101.091 101.855 101.158 ;
      RECT 101.795 98.982 101.855 101.158 ;
      RECT 99.725 101.052 101.901 101.112 ;
      RECT 101.841 98.936 101.901 101.112 ;
      RECT 99.771 101.006 101.947 101.066 ;
      RECT 101.887 98.89 101.947 101.066 ;
      RECT 99.817 100.96 101.993 101.02 ;
      RECT 101.933 98.844 101.993 101.02 ;
      RECT 99.863 100.914 102.039 100.974 ;
      RECT 101.979 98.798 102.039 100.974 ;
      RECT 99.909 100.868 102.085 100.928 ;
      RECT 102.025 98.752 102.085 100.928 ;
      RECT 99.955 100.822 102.131 100.882 ;
      RECT 102.071 98.706 102.131 100.882 ;
      RECT 100.001 100.776 102.177 100.836 ;
      RECT 102.117 98.66 102.177 100.836 ;
      RECT 100.047 100.73 102.223 100.79 ;
      RECT 102.163 98.614 102.223 100.79 ;
      RECT 100.093 100.684 102.269 100.744 ;
      RECT 102.209 98.568 102.269 100.744 ;
      RECT 100.139 100.638 102.315 100.698 ;
      RECT 102.255 98.522 102.315 100.698 ;
      RECT 100.185 100.592 102.361 100.652 ;
      RECT 102.301 98.476 102.361 100.652 ;
      RECT 100.231 100.546 102.407 100.606 ;
      RECT 102.347 98.43 102.407 100.606 ;
      RECT 100.277 100.5 102.453 100.56 ;
      RECT 102.393 98.384 102.453 100.56 ;
      RECT 102.439 98.338 102.499 100.514 ;
      RECT 102.485 98.292 102.545 100.468 ;
      RECT 102.531 98.246 102.591 100.422 ;
      RECT 102.577 98.199 102.637 100.376 ;
      RECT 102.623 98.175 102.683 100.33 ;
      RECT 102.623 98.175 102.729 100.284 ;
      RECT 102.623 98.175 102.775 100.238 ;
      RECT 102.623 98.175 102.821 100.192 ;
      RECT 102.623 98.175 102.867 100.146 ;
      RECT 102.623 98.175 102.913 100.1 ;
      RECT 102.623 98.175 102.959 100.054 ;
      RECT 102.623 98.175 103.005 100.008 ;
      RECT 102.623 98.175 103.051 99.962 ;
      RECT 102.623 98.175 103.097 99.916 ;
      RECT 102.623 98.175 103.143 99.87 ;
      RECT 102.623 98.175 103.189 99.824 ;
      RECT 102.623 98.175 103.235 99.778 ;
      RECT 102.623 98.175 103.281 99.732 ;
      RECT 102.623 98.175 103.327 99.686 ;
      RECT 102.623 98.175 103.373 99.64 ;
      RECT 102.623 98.175 103.419 99.594 ;
      RECT 102.623 98.175 103.465 99.548 ;
      RECT 102.623 98.175 103.511 99.502 ;
      RECT 102.623 98.175 103.557 99.456 ;
      RECT 102.623 98.175 103.603 99.41 ;
      RECT 102.623 98.175 103.649 99.364 ;
      RECT 101.473 99.304 103.665 99.333 ;
      RECT 102.623 98.175 110 99.325 ;
      RECT 107.675 108.902 110 110 ;
      RECT 108.925 107.675 110 110 ;
      RECT 107.721 108.856 110 110 ;
      RECT 108.917 107.679 110 110 ;
      RECT 107.767 108.81 110 110 ;
      RECT 108.871 107.706 110 110 ;
      RECT 107.813 108.764 110 110 ;
      RECT 108.825 107.752 110 110 ;
      RECT 107.859 108.718 110 110 ;
      RECT 108.779 107.798 110 110 ;
      RECT 107.905 108.672 110 110 ;
      RECT 108.733 107.844 110 110 ;
      RECT 107.951 108.626 110 110 ;
      RECT 108.687 107.89 110 110 ;
      RECT 107.997 108.58 110 110 ;
      RECT 108.641 107.936 110 110 ;
      RECT 108.043 108.534 110 110 ;
      RECT 108.595 107.982 110 110 ;
      RECT 108.089 108.488 110 110 ;
      RECT 108.549 108.028 110 110 ;
      RECT 108.135 108.442 110 110 ;
      RECT 108.503 108.074 110 110 ;
      RECT 108.181 108.396 110 110 ;
      RECT 108.457 108.12 110 110 ;
      RECT 108.227 108.35 110 110 ;
      RECT 108.411 108.166 110 110 ;
      RECT 108.273 108.304 110 110 ;
      RECT 108.365 108.212 110 110 ;
      RECT 108.319 108.258 110 110 ;
    LAYER MET5 SPACING 0.1 ;
      RECT -20 -20 3.17 110 ;
      RECT -20 -20 3.216 55.662 ;
      RECT -20 -20 3.262 55.616 ;
      RECT -20 -20 3.308 55.57 ;
      RECT -20 -20 3.354 55.524 ;
      RECT -20 -20 3.4 55.478 ;
      RECT -20 -20 3.446 55.432 ;
      RECT -20 -20 3.492 55.386 ;
      RECT -20 -20 3.538 55.34 ;
      RECT -20 -20 3.584 55.294 ;
      RECT -20 -20 3.63 55.248 ;
      RECT -20 -20 3.676 55.202 ;
      RECT -20 -20 3.722 55.156 ;
      RECT -20 -20 3.768 55.11 ;
      RECT -20 -20 3.814 55.064 ;
      RECT -20 -20 3.86 55.018 ;
      RECT -20 -20 3.906 54.972 ;
      RECT -20 -20 3.952 54.926 ;
      RECT -20 -20 3.998 54.88 ;
      RECT -20 -20 4.044 54.834 ;
      RECT -20 -20 4.09 54.788 ;
      RECT -20 -20 4.136 54.742 ;
      RECT -20 -20 4.182 54.696 ;
      RECT -20 -20 4.228 54.65 ;
      RECT -20 -20 4.274 54.604 ;
      RECT -20 -20 4.32 54.558 ;
      RECT -20 -20 4.366 54.512 ;
      RECT -20 -20 4.412 54.466 ;
      RECT -20 -20 4.458 54.42 ;
      RECT -20 -20 4.504 54.374 ;
      RECT -20 -20 4.55 54.328 ;
      RECT -20 -20 4.596 54.282 ;
      RECT -20 -20 4.642 54.236 ;
      RECT -20 -20 4.688 54.19 ;
      RECT -20 -20 4.734 54.144 ;
      RECT -20 -20 4.78 54.098 ;
      RECT -20 -20 4.826 54.052 ;
      RECT -20 -20 4.872 54.006 ;
      RECT -20 -20 4.918 53.96 ;
      RECT -20 -20 4.964 53.914 ;
      RECT -20 -20 5.01 53.868 ;
      RECT -20 -20 5.056 53.822 ;
      RECT -20 -20 5.102 53.776 ;
      RECT -20 -20 5.148 53.73 ;
      RECT -20 -20 5.194 53.684 ;
      RECT -20 -20 5.24 53.638 ;
      RECT -20 -20 5.286 53.592 ;
      RECT -20 -20 5.332 53.546 ;
      RECT -20 -20 5.378 53.5 ;
      RECT -20 -20 5.424 53.454 ;
      RECT -20 -20 5.47 53.408 ;
      RECT -20 -20 5.516 53.362 ;
      RECT -20 -20 5.562 53.316 ;
      RECT -20 -20 5.608 53.27 ;
      RECT -20 -20 5.654 53.224 ;
      RECT -20 -20 5.7 53.178 ;
      RECT -20 -20 5.746 53.132 ;
      RECT -20 -20 5.792 53.086 ;
      RECT -20 -20 5.838 53.04 ;
      RECT -20 -20 5.884 52.994 ;
      RECT -20 -20 5.93 52.948 ;
      RECT -20 -20 5.976 52.902 ;
      RECT -20 -20 6.022 52.856 ;
      RECT -20 -20 6.068 52.81 ;
      RECT -20 -20 6.114 52.764 ;
      RECT -20 -20 6.16 52.718 ;
      RECT -20 -20 6.206 52.672 ;
      RECT -20 -20 6.252 52.626 ;
      RECT -20 -20 6.298 52.58 ;
      RECT -20 -20 6.344 52.534 ;
      RECT -20 -20 6.39 52.488 ;
      RECT -20 -20 6.436 52.442 ;
      RECT -20 -20 6.482 52.396 ;
      RECT -20 -20 6.528 52.35 ;
      RECT -20 -20 6.574 52.304 ;
      RECT -20 -20 6.62 52.258 ;
      RECT -20 -20 6.666 52.212 ;
      RECT -20 -20 6.712 52.166 ;
      RECT -20 -20 6.758 52.12 ;
      RECT -20 -20 6.804 52.074 ;
      RECT -20 -20 6.85 52.028 ;
      RECT -20 -20 6.896 51.982 ;
      RECT -20 -20 6.942 51.936 ;
      RECT -20 -20 6.988 51.89 ;
      RECT -20 -20 7.034 51.844 ;
      RECT -20 -20 7.08 51.798 ;
      RECT -20 -20 7.126 51.752 ;
      RECT -20 -20 7.172 51.706 ;
      RECT -20 -20 7.218 51.66 ;
      RECT -20 -20 7.264 51.614 ;
      RECT -20 -20 7.31 51.568 ;
      RECT -20 -20 7.356 51.522 ;
      RECT -20 -20 7.402 51.476 ;
      RECT -20 -20 7.448 51.43 ;
      RECT -20 -20 7.494 51.384 ;
      RECT -20 -20 7.54 51.338 ;
      RECT -20 -20 7.586 51.292 ;
      RECT -20 -20 7.632 51.246 ;
      RECT -20 -20 7.678 51.2 ;
      RECT -20 -20 7.724 51.154 ;
      RECT -20 -20 7.77 51.108 ;
      RECT -20 -20 7.816 51.062 ;
      RECT -20 -20 7.862 51.016 ;
      RECT -20 -20 7.908 50.97 ;
      RECT -20 -20 7.954 50.924 ;
      RECT -20 -20 8 50.878 ;
      RECT -20 -20 8.046 50.832 ;
      RECT -20 -20 8.092 50.786 ;
      RECT -20 -20 8.138 50.74 ;
      RECT -20 -20 8.184 50.694 ;
      RECT -20 -20 8.23 50.648 ;
      RECT -20 -20 8.276 50.602 ;
      RECT -20 -20 8.322 50.556 ;
      RECT -20 -20 8.368 50.51 ;
      RECT -20 -20 8.414 50.464 ;
      RECT -20 -20 8.46 50.418 ;
      RECT -20 -20 8.506 50.372 ;
      RECT -20 -20 8.552 50.326 ;
      RECT -20 -20 8.598 50.28 ;
      RECT -20 -20 8.644 50.234 ;
      RECT -20 -20 8.69 50.188 ;
      RECT -20 -20 8.736 50.142 ;
      RECT -20 -20 8.782 50.096 ;
      RECT -20 -20 8.828 50.05 ;
      RECT -20 -20 8.874 50.004 ;
      RECT -20 -20 8.92 49.958 ;
      RECT -20 -20 8.966 49.912 ;
      RECT -20 -20 9.012 49.866 ;
      RECT -20 -20 9.058 49.82 ;
      RECT -20 -20 9.104 49.774 ;
      RECT -20 -20 9.15 49.728 ;
      RECT -20 -20 9.196 49.682 ;
      RECT -20 -20 9.242 49.636 ;
      RECT -20 -20 9.288 49.59 ;
      RECT -20 -20 9.334 49.544 ;
      RECT -20 -20 9.38 49.498 ;
      RECT -20 -20 9.426 49.452 ;
      RECT -20 -20 9.472 49.406 ;
      RECT -20 -20 9.518 49.36 ;
      RECT -20 -20 9.564 49.314 ;
      RECT -20 -20 9.61 49.268 ;
      RECT -20 -20 9.656 49.222 ;
      RECT -20 -20 9.702 49.176 ;
      RECT -20 -20 9.748 49.13 ;
      RECT -20 -20 9.794 49.084 ;
      RECT -20 -20 9.84 49.038 ;
      RECT -20 -20 9.886 48.992 ;
      RECT -20 -20 9.932 48.946 ;
      RECT -20 -20 9.978 48.9 ;
      RECT -20 -20 10.024 48.854 ;
      RECT -20 -20 10.07 48.808 ;
      RECT -20 -20 10.116 48.762 ;
      RECT -20 -20 10.162 48.716 ;
      RECT -20 -20 10.208 48.67 ;
      RECT -20 -20 10.254 48.624 ;
      RECT -20 -20 10.3 48.578 ;
      RECT -20 -20 10.346 48.532 ;
      RECT -20 -20 10.392 48.486 ;
      RECT -20 -20 10.438 48.44 ;
      RECT -20 -20 10.484 48.394 ;
      RECT -20 -20 10.53 48.348 ;
      RECT -20 -20 10.576 48.302 ;
      RECT -20 -20 10.622 48.256 ;
      RECT -20 -20 10.668 48.21 ;
      RECT -20 -20 10.714 48.164 ;
      RECT -20 -20 10.76 48.118 ;
      RECT -20 -20 10.806 48.072 ;
      RECT -20 -20 10.852 48.026 ;
      RECT -20 -20 10.898 47.98 ;
      RECT -20 -20 10.944 47.934 ;
      RECT -20 -20 10.99 47.888 ;
      RECT -20 -20 11.036 47.842 ;
      RECT -20 -20 11.082 47.796 ;
      RECT -20 -20 11.128 47.75 ;
      RECT -20 -20 11.174 47.704 ;
      RECT -20 -20 11.22 47.658 ;
      RECT -20 -20 11.266 47.612 ;
      RECT -20 -20 11.312 47.566 ;
      RECT -20 -20 11.358 47.52 ;
      RECT -20 -20 11.404 47.474 ;
      RECT -20 -20 11.45 47.428 ;
      RECT -20 -20 11.496 47.382 ;
      RECT -20 -20 11.542 47.336 ;
      RECT -20 -20 11.588 47.29 ;
      RECT -20 -20 11.634 47.244 ;
      RECT -20 -20 11.68 47.198 ;
      RECT -20 -20 11.726 47.152 ;
      RECT -20 -20 11.772 47.106 ;
      RECT -20 -20 11.818 47.06 ;
      RECT -20 -20 11.864 47.014 ;
      RECT -20 -20 11.91 46.968 ;
      RECT -20 -20 11.956 46.922 ;
      RECT -20 -20 12.002 46.876 ;
      RECT -20 -20 12.048 46.83 ;
      RECT -20 -20 12.094 46.784 ;
      RECT -20 -20 12.14 46.738 ;
      RECT -20 -20 12.186 46.692 ;
      RECT -20 -20 12.232 46.646 ;
      RECT -20 -20 12.278 46.6 ;
      RECT -20 -20 12.324 46.554 ;
      RECT -20 -20 12.37 46.508 ;
      RECT -20 -20 12.416 46.462 ;
      RECT -20 -20 12.462 46.416 ;
      RECT -20 -20 12.508 46.37 ;
      RECT -20 -20 12.554 46.324 ;
      RECT -20 -20 12.6 46.278 ;
      RECT -20 -20 12.646 46.232 ;
      RECT -20 -20 12.692 46.186 ;
      RECT -20 -20 12.738 46.14 ;
      RECT -20 -20 12.784 46.094 ;
      RECT -20 -20 12.83 46.048 ;
      RECT -20 -20 12.876 46.002 ;
      RECT -20 -20 12.922 45.956 ;
      RECT -20 -20 12.968 45.91 ;
      RECT -20 -20 13.014 45.864 ;
      RECT -20 -20 13.06 45.818 ;
      RECT -20 -20 13.106 45.772 ;
      RECT -20 -20 13.152 45.726 ;
      RECT -20 -20 13.198 45.68 ;
      RECT -20 -20 13.244 45.634 ;
      RECT -20 -20 13.29 45.588 ;
      RECT -20 -20 13.336 45.542 ;
      RECT -20 -20 13.382 45.496 ;
      RECT -20 -20 13.428 45.45 ;
      RECT -20 -20 13.474 45.404 ;
      RECT -20 -20 13.52 45.358 ;
      RECT -20 -20 13.566 45.312 ;
      RECT -20 -20 13.612 45.266 ;
      RECT -20 -20 13.658 45.22 ;
      RECT -20 -20 13.704 45.174 ;
      RECT -20 -20 13.75 45.128 ;
      RECT -20 -20 13.796 45.082 ;
      RECT -20 -20 13.842 45.036 ;
      RECT -20 -20 13.888 44.99 ;
      RECT -20 -20 13.934 44.944 ;
      RECT -20 -20 13.98 44.898 ;
      RECT -20 -20 14.026 44.852 ;
      RECT -20 -20 14.072 44.806 ;
      RECT -20 -20 14.118 44.76 ;
      RECT -20 -20 14.164 44.714 ;
      RECT -20 -20 14.21 44.668 ;
      RECT -20 -20 14.256 44.622 ;
      RECT -20 -20 14.302 44.576 ;
      RECT -20 -20 14.348 44.53 ;
      RECT -20 -20 14.394 44.484 ;
      RECT -20 -20 14.44 44.438 ;
      RECT -20 -20 14.486 44.392 ;
      RECT -20 -20 14.532 44.346 ;
      RECT -20 -20 14.578 44.3 ;
      RECT -20 -20 14.624 44.254 ;
      RECT -20 -20 14.67 44.208 ;
      RECT -20 -20 14.716 44.162 ;
      RECT -20 -20 14.762 44.116 ;
      RECT -20 -20 14.808 44.07 ;
      RECT -20 -20 14.854 44.024 ;
      RECT -20 -20 14.9 43.978 ;
      RECT -20 -20 14.946 43.932 ;
      RECT -20 -20 14.992 43.886 ;
      RECT -20 -20 15.038 43.84 ;
      RECT -20 -20 15.084 43.794 ;
      RECT -20 -20 15.13 43.748 ;
      RECT -20 -20 15.17 43.705 ;
      RECT -20 -20 15.216 43.662 ;
      RECT -20 -20 15.262 43.616 ;
      RECT -20 -20 15.308 43.57 ;
      RECT -20 -20 15.354 43.524 ;
      RECT -20 -20 15.4 43.478 ;
      RECT -20 -20 15.446 43.432 ;
      RECT -20 -20 15.492 43.386 ;
      RECT -20 -20 15.538 43.34 ;
      RECT -20 -20 15.584 43.294 ;
      RECT -20 -20 15.63 43.248 ;
      RECT -20 -20 15.676 43.202 ;
      RECT -20 -20 15.722 43.156 ;
      RECT -20 -20 15.768 43.11 ;
      RECT -20 -20 15.814 43.064 ;
      RECT -20 -20 15.86 43.018 ;
      RECT -20 -20 15.906 42.972 ;
      RECT -20 -20 15.952 42.926 ;
      RECT -20 -20 15.998 42.88 ;
      RECT -20 -20 16.044 42.834 ;
      RECT -20 -20 16.09 42.788 ;
      RECT -20 -20 16.136 42.742 ;
      RECT -20 -20 16.182 42.696 ;
      RECT -20 -20 16.228 42.65 ;
      RECT -20 -20 16.274 42.604 ;
      RECT -20 -20 16.32 42.558 ;
      RECT -20 -20 16.366 42.512 ;
      RECT -20 -20 16.412 42.466 ;
      RECT -20 -20 16.458 42.42 ;
      RECT -20 -20 16.504 42.374 ;
      RECT -20 -20 16.55 42.328 ;
      RECT -20 -20 16.596 42.282 ;
      RECT -20 -20 16.642 42.236 ;
      RECT -20 -20 16.688 42.19 ;
      RECT -20 -20 16.734 42.144 ;
      RECT -20 -20 16.78 42.098 ;
      RECT -20 -20 16.826 42.052 ;
      RECT -20 -20 16.872 42.006 ;
      RECT -20 -20 16.918 41.96 ;
      RECT -20 -20 16.964 41.914 ;
      RECT -20 -20 17.01 41.868 ;
      RECT -20 -20 17.056 41.822 ;
      RECT -20 -20 17.102 41.776 ;
      RECT -20 -20 17.148 41.73 ;
      RECT -20 -20 17.194 41.684 ;
      RECT -20 -20 17.24 41.638 ;
      RECT -20 -20 17.286 41.592 ;
      RECT -20 -20 17.332 41.546 ;
      RECT -20 -20 17.378 41.5 ;
      RECT -20 -20 17.424 41.454 ;
      RECT -20 -20 17.47 41.408 ;
      RECT -20 -20 17.516 41.362 ;
      RECT -20 -20 17.562 41.316 ;
      RECT -20 -20 17.608 41.27 ;
      RECT -20 -20 17.654 41.224 ;
      RECT -20 -20 17.7 41.178 ;
      RECT -20 -20 17.746 41.132 ;
      RECT -20 -20 17.792 41.086 ;
      RECT -20 -20 17.838 41.04 ;
      RECT -20 -20 17.884 40.994 ;
      RECT -20 -20 17.93 40.948 ;
      RECT -20 -20 17.976 40.902 ;
      RECT -20 -20 18.022 40.856 ;
      RECT -20 -20 18.068 40.81 ;
      RECT -20 -20 18.114 40.764 ;
      RECT -20 -20 18.16 40.718 ;
      RECT -20 -20 18.206 40.672 ;
      RECT -20 -20 18.252 40.626 ;
      RECT -20 -20 18.298 40.58 ;
      RECT -20 -20 18.344 40.534 ;
      RECT -20 -20 18.39 40.488 ;
      RECT -20 -20 18.436 40.442 ;
      RECT -20 -20 18.482 40.396 ;
      RECT -20 -20 18.528 40.35 ;
      RECT -20 -20 18.574 40.304 ;
      RECT -20 -20 18.62 40.258 ;
      RECT -20 -20 18.666 40.212 ;
      RECT -20 -20 18.712 40.166 ;
      RECT -20 -20 18.758 40.12 ;
      RECT -20 -20 18.804 40.074 ;
      RECT -20 -20 18.85 40.028 ;
      RECT -20 -20 18.896 39.982 ;
      RECT -20 -20 18.942 39.936 ;
      RECT -20 -20 18.988 39.89 ;
      RECT -20 -20 19.034 39.844 ;
      RECT -20 -20 19.08 39.798 ;
      RECT -20 -20 19.126 39.752 ;
      RECT -20 -20 19.172 39.706 ;
      RECT -20 -20 19.218 39.66 ;
      RECT -20 -20 19.264 39.614 ;
      RECT -20 -20 19.31 39.568 ;
      RECT -20 -20 19.356 39.522 ;
      RECT -20 -20 19.402 39.476 ;
      RECT -20 -20 19.448 39.43 ;
      RECT -20 -20 19.494 39.384 ;
      RECT -20 -20 19.54 39.338 ;
      RECT -20 -20 19.586 39.292 ;
      RECT -20 -20 19.632 39.246 ;
      RECT -20 -20 19.678 39.2 ;
      RECT -20 -20 19.724 39.154 ;
      RECT -20 -20 19.77 39.108 ;
      RECT -20 -20 19.816 39.062 ;
      RECT -20 -20 19.862 39.016 ;
      RECT -20 -20 19.908 38.97 ;
      RECT -20 -20 19.954 38.924 ;
      RECT -20 -20 20 38.878 ;
      RECT -20 -20 20.046 38.832 ;
      RECT -20 -20 20.092 38.786 ;
      RECT -20 -20 20.138 38.74 ;
      RECT -20 -20 20.184 38.694 ;
      RECT -20 -20 20.23 38.648 ;
      RECT -20 -20 20.276 38.602 ;
      RECT -20 -20 20.322 38.556 ;
      RECT -20 -20 20.368 38.51 ;
      RECT -20 -20 20.414 38.464 ;
      RECT -20 -20 20.46 38.418 ;
      RECT -20 -20 20.506 38.372 ;
      RECT -20 -20 20.552 38.326 ;
      RECT -20 -20 20.598 38.28 ;
      RECT -20 -20 20.644 38.234 ;
      RECT -20 -20 20.69 38.188 ;
      RECT -20 -20 20.736 38.142 ;
      RECT -20 -20 20.782 38.096 ;
      RECT -20 -20 20.828 38.05 ;
      RECT -20 -20 20.874 38.004 ;
      RECT -20 -20 20.92 37.958 ;
      RECT -20 -20 20.966 37.912 ;
      RECT -20 -20 21.012 37.866 ;
      RECT -20 -20 21.058 37.82 ;
      RECT -20 -20 21.104 37.774 ;
      RECT -20 -20 21.15 37.728 ;
      RECT -20 -20 21.196 37.682 ;
      RECT -20 -20 21.242 37.636 ;
      RECT -20 -20 21.288 37.59 ;
      RECT -20 -20 21.334 37.544 ;
      RECT -20 -20 21.38 37.498 ;
      RECT -20 -20 21.426 37.452 ;
      RECT -20 -20 21.472 37.406 ;
      RECT -20 -20 21.518 37.36 ;
      RECT -20 -20 21.564 37.314 ;
      RECT -20 -20 21.61 37.268 ;
      RECT -20 -20 21.656 37.222 ;
      RECT -20 -20 21.702 37.176 ;
      RECT -20 -20 21.748 37.13 ;
      RECT -20 -20 21.794 37.084 ;
      RECT -20 -20 21.84 37.038 ;
      RECT -20 -20 21.886 36.992 ;
      RECT -20 -20 21.932 36.946 ;
      RECT -20 -20 21.978 36.9 ;
      RECT -20 -20 22.024 36.854 ;
      RECT -20 -20 22.07 36.808 ;
      RECT -20 -20 22.116 36.762 ;
      RECT -20 -20 22.162 36.716 ;
      RECT -20 -20 22.208 36.67 ;
      RECT -20 -20 22.254 36.624 ;
      RECT -20 -20 22.3 36.578 ;
      RECT -20 -20 22.346 36.532 ;
      RECT -20 -20 22.392 36.486 ;
      RECT -20 -20 22.438 36.44 ;
      RECT -20 -20 22.484 36.394 ;
      RECT -20 -20 22.53 36.348 ;
      RECT -20 -20 22.576 36.302 ;
      RECT -20 -20 22.622 36.256 ;
      RECT -20 -20 22.668 36.21 ;
      RECT -20 -20 22.714 36.164 ;
      RECT -20 -20 22.76 36.118 ;
      RECT -20 -20 22.806 36.072 ;
      RECT -20 -20 22.852 36.026 ;
      RECT -20 -20 22.898 35.98 ;
      RECT -20 -20 22.944 35.934 ;
      RECT -20 -20 22.99 35.888 ;
      RECT -20 -20 23.036 35.842 ;
      RECT -20 -20 23.082 35.796 ;
      RECT -20 -20 23.128 35.75 ;
      RECT -20 -20 23.174 35.704 ;
      RECT -20 -20 23.22 35.658 ;
      RECT -20 -20 23.266 35.612 ;
      RECT -20 -20 23.312 35.566 ;
      RECT -20 -20 23.358 35.52 ;
      RECT -20 -20 23.404 35.474 ;
      RECT -20 -20 23.45 35.428 ;
      RECT -20 -20 23.496 35.382 ;
      RECT -20 -20 23.542 35.336 ;
      RECT -20 -20 23.588 35.29 ;
      RECT -20 -20 23.634 35.244 ;
      RECT -20 -20 23.68 35.198 ;
      RECT -20 -20 23.726 35.152 ;
      RECT -20 -20 23.772 35.106 ;
      RECT -20 -20 23.818 35.06 ;
      RECT -20 -20 23.864 35.014 ;
      RECT -20 -20 23.91 34.968 ;
      RECT -20 -20 23.956 34.922 ;
      RECT -20 -20 24.002 34.876 ;
      RECT -20 -20 24.048 34.83 ;
      RECT -20 -20 24.094 34.784 ;
      RECT -20 -20 24.14 34.738 ;
      RECT -20 -20 24.186 34.692 ;
      RECT -20 -20 24.232 34.646 ;
      RECT -20 -20 24.278 34.6 ;
      RECT -20 -20 24.324 34.554 ;
      RECT -20 -20 24.37 34.508 ;
      RECT -20 -20 24.416 34.462 ;
      RECT -20 -20 24.462 34.416 ;
      RECT -20 -20 24.508 34.37 ;
      RECT -20 -20 24.554 34.324 ;
      RECT -20 -20 24.6 34.278 ;
      RECT -20 -20 24.646 34.232 ;
      RECT -20 -20 24.692 34.186 ;
      RECT -20 -20 24.738 34.14 ;
      RECT -20 -20 24.784 34.094 ;
      RECT -20 -20 24.83 34.048 ;
      RECT -20 -20 24.876 34.002 ;
      RECT -20 -20 24.922 33.956 ;
      RECT -20 -20 24.968 33.91 ;
      RECT -20 -20 25.014 33.864 ;
      RECT -20 -20 25.06 33.818 ;
      RECT -20 -20 25.106 33.772 ;
      RECT -20 -20 25.152 33.726 ;
      RECT -20 -20 25.198 33.68 ;
      RECT -20 -20 25.244 33.634 ;
      RECT -20 -20 25.29 33.588 ;
      RECT -20 -20 25.336 33.542 ;
      RECT -20 -20 25.382 33.496 ;
      RECT -20 -20 25.428 33.45 ;
      RECT -20 -20 25.474 33.404 ;
      RECT -20 -20 25.52 33.358 ;
      RECT -20 -20 25.566 33.312 ;
      RECT -20 -20 25.612 33.266 ;
      RECT -20 -20 25.658 33.22 ;
      RECT -20 -20 25.704 33.174 ;
      RECT -20 -20 25.75 33.128 ;
      RECT -20 -20 25.796 33.082 ;
      RECT -20 -20 25.842 33.036 ;
      RECT -20 -20 25.888 32.99 ;
      RECT -20 -20 25.934 32.944 ;
      RECT -20 -20 25.98 32.898 ;
      RECT -20 -20 26.026 32.852 ;
      RECT -20 -20 26.072 32.806 ;
      RECT -20 -20 26.118 32.76 ;
      RECT -20 -20 26.164 32.714 ;
      RECT -20 -20 26.21 32.668 ;
      RECT -20 -20 26.256 32.622 ;
      RECT -20 -20 26.302 32.576 ;
      RECT -20 -20 26.348 32.53 ;
      RECT -20 -20 26.394 32.484 ;
      RECT -20 -20 26.44 32.438 ;
      RECT -20 -20 26.486 32.392 ;
      RECT -20 -20 26.532 32.346 ;
      RECT -20 -20 26.578 32.3 ;
      RECT -20 -20 26.624 32.254 ;
      RECT -20 -20 26.67 32.208 ;
      RECT -20 -20 26.716 32.162 ;
      RECT -20 -20 26.762 32.116 ;
      RECT -20 -20 26.808 32.07 ;
      RECT -20 -20 26.854 32.024 ;
      RECT -20 -20 26.9 31.978 ;
      RECT -20 -20 26.946 31.932 ;
      RECT -20 -20 26.992 31.886 ;
      RECT -20 -20 27.038 31.84 ;
      RECT -20 -20 27.084 31.794 ;
      RECT -20 -20 27.13 31.748 ;
      RECT -20 -20 27.176 31.702 ;
      RECT -20 -20 27.222 31.656 ;
      RECT -20 -20 27.268 31.61 ;
      RECT -20 -20 27.314 31.564 ;
      RECT -20 -20 27.36 31.518 ;
      RECT -20 -20 27.406 31.472 ;
      RECT -20 -20 27.452 31.426 ;
      RECT -20 -20 27.498 31.38 ;
      RECT -20 -20 27.544 31.334 ;
      RECT -20 -20 27.59 31.288 ;
      RECT -20 -20 27.636 31.242 ;
      RECT -20 -20 27.682 31.196 ;
      RECT -20 -20 27.728 31.15 ;
      RECT -20 -20 27.774 31.104 ;
      RECT -20 -20 27.82 31.058 ;
      RECT -20 -20 27.866 31.012 ;
      RECT -20 -20 27.912 30.966 ;
      RECT -20 -20 27.958 30.92 ;
      RECT -20 -20 28.004 30.874 ;
      RECT -20 -20 28.05 30.828 ;
      RECT -20 -20 28.096 30.782 ;
      RECT -20 -20 28.142 30.736 ;
      RECT -20 -20 28.188 30.69 ;
      RECT -20 -20 28.234 30.644 ;
      RECT -20 -20 28.28 30.598 ;
      RECT -20 -20 28.326 30.552 ;
      RECT -20 -20 28.372 30.506 ;
      RECT -20 -20 28.418 30.46 ;
      RECT -20 -20 28.464 30.414 ;
      RECT -20 -20 28.51 30.368 ;
      RECT -20 -20 28.556 30.322 ;
      RECT -20 -20 28.602 30.276 ;
      RECT -20 -20 28.648 30.23 ;
      RECT -20 -20 28.694 30.184 ;
      RECT -20 -20 28.74 30.138 ;
      RECT -20 -20 28.786 30.092 ;
      RECT -20 -20 28.832 30.046 ;
      RECT -20 -20 28.878 30 ;
      RECT -20 -20 28.924 29.954 ;
      RECT -20 -20 28.97 29.908 ;
      RECT -20 -20 29.016 29.862 ;
      RECT -20 -20 29.062 29.816 ;
      RECT -20 -20 29.108 29.77 ;
      RECT -20 -20 29.154 29.724 ;
      RECT -20 -20 29.2 29.678 ;
      RECT -20 -20 29.246 29.632 ;
      RECT -20 -20 29.292 29.586 ;
      RECT -20 -20 29.338 29.54 ;
      RECT -20 -20 29.384 29.494 ;
      RECT -20 -20 29.43 29.448 ;
      RECT -20 -20 29.476 29.402 ;
      RECT -20 -20 29.522 29.356 ;
      RECT -20 -20 29.568 29.31 ;
      RECT -20 -20 29.614 29.264 ;
      RECT -20 -20 29.66 29.218 ;
      RECT -20 -20 29.706 29.172 ;
      RECT -20 -20 29.752 29.126 ;
      RECT -20 -20 29.798 29.08 ;
      RECT -20 -20 29.844 29.034 ;
      RECT -20 -20 29.89 28.988 ;
      RECT -20 -20 29.936 28.942 ;
      RECT -20 -20 29.982 28.896 ;
      RECT -20 -20 30.028 28.85 ;
      RECT -20 -20 30.074 28.804 ;
      RECT -20 -20 30.12 28.758 ;
      RECT -20 -20 30.166 28.712 ;
      RECT -20 -20 30.212 28.666 ;
      RECT -20 -20 30.258 28.62 ;
      RECT -20 -20 30.304 28.574 ;
      RECT -20 -20 30.35 28.528 ;
      RECT -20 -20 30.396 28.482 ;
      RECT -20 -20 30.442 28.436 ;
      RECT -20 -20 30.488 28.39 ;
      RECT -20 -20 30.534 28.344 ;
      RECT -20 -20 30.58 28.298 ;
      RECT -20 -20 30.626 28.252 ;
      RECT -20 -20 30.672 28.206 ;
      RECT -20 -20 30.718 28.16 ;
      RECT -20 -20 30.764 28.114 ;
      RECT -20 -20 30.81 28.068 ;
      RECT -20 -20 30.856 28.022 ;
      RECT -20 -20 30.902 27.976 ;
      RECT -20 -20 30.948 27.93 ;
      RECT -20 -20 30.994 27.884 ;
      RECT -20 -20 31.04 27.838 ;
      RECT -20 -20 31.086 27.792 ;
      RECT -20 -20 31.132 27.746 ;
      RECT -20 -20 31.178 27.7 ;
      RECT -20 -20 31.224 27.654 ;
      RECT -20 -20 31.27 27.608 ;
      RECT -20 -20 31.316 27.562 ;
      RECT -20 -20 31.362 27.516 ;
      RECT -20 -20 31.408 27.47 ;
      RECT -20 -20 31.454 27.424 ;
      RECT -20 -20 31.5 27.378 ;
      RECT -20 -20 31.546 27.332 ;
      RECT -20 -20 31.592 27.286 ;
      RECT -20 -20 31.638 27.24 ;
      RECT -20 -20 31.684 27.194 ;
      RECT -20 -20 31.73 27.148 ;
      RECT -20 -20 31.776 27.102 ;
      RECT -20 -20 31.822 27.056 ;
      RECT -20 -20 31.868 27.01 ;
      RECT -20 -20 31.914 26.964 ;
      RECT -20 -20 31.96 26.918 ;
      RECT -20 -20 32.006 26.872 ;
      RECT -20 -20 32.052 26.826 ;
      RECT -20 -20 32.098 26.78 ;
      RECT -20 -20 32.144 26.734 ;
      RECT -20 -20 32.19 26.688 ;
      RECT -20 -20 32.236 26.642 ;
      RECT -20 -20 32.282 26.596 ;
      RECT -20 -20 32.328 26.55 ;
      RECT -20 -20 32.374 26.504 ;
      RECT -20 -20 32.42 26.458 ;
      RECT -20 -20 32.466 26.412 ;
      RECT -20 -20 32.512 26.366 ;
      RECT -20 -20 32.558 26.32 ;
      RECT -20 -20 32.604 26.274 ;
      RECT -20 -20 32.65 26.228 ;
      RECT -20 -20 32.696 26.182 ;
      RECT -20 -20 32.742 26.136 ;
      RECT -20 -20 32.788 26.09 ;
      RECT -20 -20 32.834 26.044 ;
      RECT -20 -20 32.88 25.998 ;
      RECT -20 -20 32.926 25.952 ;
      RECT -20 -20 32.972 25.906 ;
      RECT -20 -20 33.018 25.86 ;
      RECT -20 -20 33.064 25.814 ;
      RECT -20 -20 33.11 25.768 ;
      RECT -20 -20 33.156 25.722 ;
      RECT -20 -20 33.202 25.676 ;
      RECT -20 -20 33.248 25.63 ;
      RECT -20 -20 33.294 25.584 ;
      RECT -20 -20 33.34 25.538 ;
      RECT -20 -20 33.386 25.492 ;
      RECT -20 -20 33.432 25.446 ;
      RECT -20 -20 33.478 25.4 ;
      RECT -20 -20 33.524 25.354 ;
      RECT -20 -20 33.57 25.308 ;
      RECT -20 -20 33.616 25.262 ;
      RECT -20 -20 33.662 25.216 ;
      RECT -20 -20 33.708 25.17 ;
      RECT -20 -20 33.754 25.124 ;
      RECT -20 -20 33.8 25.078 ;
      RECT -20 -20 33.846 25.032 ;
      RECT -20 -20 33.892 24.986 ;
      RECT -20 -20 33.938 24.94 ;
      RECT -20 -20 33.984 24.894 ;
      RECT -20 -20 34.03 24.848 ;
      RECT -20 -20 34.076 24.802 ;
      RECT -20 -20 34.122 24.756 ;
      RECT -20 -20 34.168 24.71 ;
      RECT -20 -20 34.214 24.664 ;
      RECT -20 -20 34.26 24.618 ;
      RECT -20 -20 34.306 24.572 ;
      RECT -20 -20 34.352 24.526 ;
      RECT -20 -20 34.398 24.48 ;
      RECT -20 -20 34.444 24.434 ;
      RECT -20 -20 34.49 24.388 ;
      RECT -20 -20 34.536 24.342 ;
      RECT -20 -20 34.582 24.296 ;
      RECT -20 -20 34.628 24.25 ;
      RECT -20 -20 34.674 24.204 ;
      RECT -20 -20 34.72 24.158 ;
      RECT -20 -20 34.766 24.112 ;
      RECT -20 -20 34.812 24.066 ;
      RECT -20 -20 34.858 24.02 ;
      RECT -20 -20 34.904 23.974 ;
      RECT -20 -20 34.95 23.928 ;
      RECT -20 -20 34.996 23.882 ;
      RECT -20 -20 35.042 23.836 ;
      RECT -20 -20 35.088 23.79 ;
      RECT -20 -20 35.134 23.744 ;
      RECT -20 -20 35.18 23.698 ;
      RECT -20 -20 35.226 23.652 ;
      RECT -20 -20 35.272 23.606 ;
      RECT -20 -20 35.318 23.56 ;
      RECT -20 -20 35.364 23.514 ;
      RECT -20 -20 35.41 23.468 ;
      RECT -20 -20 35.456 23.422 ;
      RECT -20 -20 35.502 23.376 ;
      RECT -20 -20 35.548 23.33 ;
      RECT -20 -20 35.594 23.284 ;
      RECT -20 -20 35.64 23.238 ;
      RECT -20 -20 35.686 23.192 ;
      RECT -20 -20 35.732 23.146 ;
      RECT -20 -20 35.778 23.1 ;
      RECT -20 -20 35.824 23.054 ;
      RECT -20 -20 35.87 23.008 ;
      RECT -20 -20 35.916 22.962 ;
      RECT -20 -20 35.962 22.916 ;
      RECT -20 -20 36.008 22.87 ;
      RECT -20 -20 36.054 22.824 ;
      RECT -20 -20 36.1 22.778 ;
      RECT -20 -20 36.146 22.732 ;
      RECT -20 -20 36.192 22.686 ;
      RECT -20 -20 36.238 22.64 ;
      RECT -20 -20 36.284 22.594 ;
      RECT -20 -20 36.33 22.548 ;
      RECT -20 -20 36.376 22.502 ;
      RECT -20 -20 36.422 22.456 ;
      RECT -20 -20 36.468 22.41 ;
      RECT -20 -20 36.514 22.364 ;
      RECT -20 -20 36.56 22.318 ;
      RECT -20 -20 36.606 22.272 ;
      RECT -20 -20 36.652 22.226 ;
      RECT -20 -20 36.698 22.18 ;
      RECT -20 -20 36.744 22.134 ;
      RECT -20 -20 36.79 22.088 ;
      RECT -20 -20 36.836 22.042 ;
      RECT -20 -20 36.882 21.996 ;
      RECT -20 -20 36.928 21.95 ;
      RECT -20 -20 36.974 21.904 ;
      RECT -20 -20 37.02 21.858 ;
      RECT -20 -20 37.066 21.812 ;
      RECT -20 -20 37.112 21.766 ;
      RECT -20 -20 37.158 21.72 ;
      RECT -20 -20 37.204 21.674 ;
      RECT -20 -20 37.25 21.628 ;
      RECT -20 -20 37.296 21.582 ;
      RECT -20 -20 37.342 21.536 ;
      RECT -20 -20 37.388 21.49 ;
      RECT -20 -20 37.434 21.444 ;
      RECT -20 -20 37.48 21.398 ;
      RECT -20 -20 37.526 21.352 ;
      RECT -20 -20 37.572 21.306 ;
      RECT -20 -20 37.618 21.26 ;
      RECT -20 -20 37.664 21.214 ;
      RECT -20 -20 37.71 21.168 ;
      RECT -20 -20 37.756 21.122 ;
      RECT -20 -20 37.802 21.076 ;
      RECT -20 -20 37.848 21.03 ;
      RECT -20 -20 37.894 20.984 ;
      RECT -20 -20 37.94 20.938 ;
      RECT -20 -20 37.986 20.892 ;
      RECT -20 -20 38.032 20.846 ;
      RECT -20 -20 38.078 20.8 ;
      RECT -20 -20 38.124 20.754 ;
      RECT -20 -20 38.17 20.708 ;
      RECT -20 -20 38.216 20.662 ;
      RECT -20 -20 38.262 20.616 ;
      RECT -20 -20 38.308 20.57 ;
      RECT -20 -20 38.354 20.524 ;
      RECT -20 -20 38.4 20.478 ;
      RECT -20 -20 38.446 20.432 ;
      RECT -20 -20 38.492 20.386 ;
      RECT -20 -20 38.538 20.34 ;
      RECT -20 -20 38.584 20.294 ;
      RECT -20 -20 38.63 20.248 ;
      RECT -20 -20 38.676 20.202 ;
      RECT -20 -20 38.722 20.156 ;
      RECT -20 -20 38.768 20.11 ;
      RECT -20 -20 38.814 20.064 ;
      RECT -20 -20 38.86 20.018 ;
      RECT -20 -20 38.906 19.972 ;
      RECT -20 -20 38.952 19.926 ;
      RECT -20 -20 38.998 19.88 ;
      RECT -20 -20 39.044 19.834 ;
      RECT -20 -20 39.09 19.788 ;
      RECT -20 -20 39.136 19.742 ;
      RECT -20 -20 39.182 19.696 ;
      RECT -20 -20 39.228 19.65 ;
      RECT -20 -20 39.274 19.604 ;
      RECT -20 -20 39.32 19.558 ;
      RECT -20 -20 39.366 19.512 ;
      RECT -20 -20 39.412 19.466 ;
      RECT -20 -20 39.458 19.42 ;
      RECT -20 -20 39.504 19.374 ;
      RECT -20 -20 39.55 19.328 ;
      RECT -20 -20 39.596 19.282 ;
      RECT -20 -20 39.642 19.236 ;
      RECT -20 -20 39.688 19.19 ;
      RECT -20 -20 39.734 19.144 ;
      RECT -20 -20 39.78 19.098 ;
      RECT -20 -20 39.826 19.052 ;
      RECT -20 -20 39.872 19.006 ;
      RECT -20 -20 39.918 18.96 ;
      RECT -20 -20 39.964 18.914 ;
      RECT -20 -20 40.01 18.868 ;
      RECT -20 -20 40.056 18.822 ;
      RECT -20 -20 40.102 18.776 ;
      RECT -20 -20 40.148 18.73 ;
      RECT -20 -20 40.194 18.684 ;
      RECT -20 -20 40.24 18.638 ;
      RECT -20 -20 40.286 18.592 ;
      RECT -20 -20 40.332 18.546 ;
      RECT -20 -20 40.378 18.5 ;
      RECT -20 -20 40.424 18.454 ;
      RECT -20 -20 40.47 18.408 ;
      RECT -20 -20 40.516 18.362 ;
      RECT -20 -20 40.562 18.316 ;
      RECT -20 -20 40.608 18.27 ;
      RECT -20 -20 40.654 18.224 ;
      RECT -20 -20 40.7 18.178 ;
      RECT -20 -20 40.746 18.132 ;
      RECT -20 -20 40.792 18.086 ;
      RECT -20 -20 40.838 18.04 ;
      RECT -20 -20 40.884 17.994 ;
      RECT -20 -20 40.93 17.948 ;
      RECT -20 -20 40.976 17.902 ;
      RECT -20 -20 41.022 17.856 ;
      RECT -20 -20 41.068 17.81 ;
      RECT -20 -20 41.114 17.764 ;
      RECT -20 -20 41.16 17.718 ;
      RECT -20 -20 41.206 17.672 ;
      RECT -20 -20 41.252 17.626 ;
      RECT -20 -20 41.298 17.58 ;
      RECT -20 -20 41.344 17.534 ;
      RECT -20 -20 41.39 17.488 ;
      RECT -20 -20 41.436 17.442 ;
      RECT -20 -20 41.482 17.396 ;
      RECT -20 -20 41.528 17.35 ;
      RECT -20 -20 41.574 17.304 ;
      RECT -20 -20 41.62 17.258 ;
      RECT -20 -20 41.666 17.212 ;
      RECT -20 -20 41.712 17.166 ;
      RECT -20 -20 41.758 17.12 ;
      RECT -20 -20 41.804 17.074 ;
      RECT -20 -20 41.85 17.028 ;
      RECT -20 -20 41.896 16.982 ;
      RECT -20 -20 41.942 16.936 ;
      RECT -20 -20 41.988 16.89 ;
      RECT -20 -20 42.034 16.844 ;
      RECT -20 -20 42.08 16.798 ;
      RECT -20 -20 42.126 16.752 ;
      RECT -20 -20 42.172 16.706 ;
      RECT -20 -20 42.218 16.66 ;
      RECT -20 -20 42.264 16.614 ;
      RECT -20 -20 42.31 16.568 ;
      RECT -20 -20 42.356 16.522 ;
      RECT -20 -20 42.402 16.476 ;
      RECT -20 -20 42.448 16.43 ;
      RECT -20 -20 42.494 16.384 ;
      RECT -20 -20 42.54 16.338 ;
      RECT -20 -20 42.586 16.292 ;
      RECT -20 -20 42.632 16.246 ;
      RECT -20 -20 42.678 16.2 ;
      RECT -20 -20 42.724 16.154 ;
      RECT -20 -20 42.77 16.108 ;
      RECT -20 -20 42.816 16.062 ;
      RECT -20 -20 42.862 16.016 ;
      RECT -20 -20 42.908 15.97 ;
      RECT -20 -20 42.954 15.924 ;
      RECT -20 -20 43 15.878 ;
      RECT -20 -20 43.046 15.832 ;
      RECT -20 -20 43.092 15.786 ;
      RECT -20 -20 43.138 15.74 ;
      RECT -20 -20 43.184 15.694 ;
      RECT -20 -20 43.23 15.648 ;
      RECT -20 -20 43.276 15.602 ;
      RECT -20 -20 43.322 15.556 ;
      RECT -20 -20 43.368 15.51 ;
      RECT -20 -20 43.414 15.464 ;
      RECT -20 -20 43.46 15.418 ;
      RECT -20 -20 43.506 15.372 ;
      RECT -20 -20 43.552 15.326 ;
      RECT -20 -20 43.598 15.28 ;
      RECT -20 -20 43.644 15.234 ;
      RECT -20 -20 43.69 15.188 ;
      RECT -20 -20 43.736 15.142 ;
      RECT -20 -20 43.782 15.096 ;
      RECT -20 -20 43.828 15.05 ;
      RECT -20 -20 43.874 15.004 ;
      RECT -20 -20 43.92 14.958 ;
      RECT -20 -20 43.966 14.912 ;
      RECT -20 -20 44.012 14.866 ;
      RECT -20 -20 44.058 14.82 ;
      RECT -20 -20 44.104 14.774 ;
      RECT -20 -20 44.15 14.728 ;
      RECT -20 -20 44.196 14.682 ;
      RECT -20 -20 44.242 14.636 ;
      RECT -20 -20 44.288 14.59 ;
      RECT -20 -20 44.334 14.544 ;
      RECT -20 -20 44.38 14.498 ;
      RECT -20 -20 44.426 14.452 ;
      RECT -20 -20 44.472 14.406 ;
      RECT -20 -20 44.518 14.36 ;
      RECT -20 -20 44.564 14.314 ;
      RECT -20 -20 44.61 14.268 ;
      RECT -20 -20 44.656 14.222 ;
      RECT -20 -20 44.702 14.176 ;
      RECT -20 -20 44.748 14.13 ;
      RECT -20 -20 44.794 14.084 ;
      RECT -20 -20 44.84 14.038 ;
      RECT -20 -20 44.886 13.992 ;
      RECT -20 -20 44.932 13.946 ;
      RECT -20 -20 44.978 13.9 ;
      RECT -20 -20 45.024 13.854 ;
      RECT -20 -20 45.07 13.808 ;
      RECT -20 -20 45.116 13.762 ;
      RECT -20 -20 45.162 13.716 ;
      RECT -20 -20 45.208 13.67 ;
      RECT -20 -20 45.254 13.624 ;
      RECT -20 -20 45.3 13.578 ;
      RECT -20 -20 45.346 13.532 ;
      RECT -20 -20 45.392 13.486 ;
      RECT -20 -20 45.438 13.44 ;
      RECT -20 -20 45.484 13.394 ;
      RECT -20 -20 45.53 13.348 ;
      RECT -20 -20 45.576 13.302 ;
      RECT -20 -20 45.622 13.256 ;
      RECT -20 -20 45.668 13.21 ;
      RECT -20 -20 45.714 13.164 ;
      RECT -20 -20 45.76 13.118 ;
      RECT -20 -20 45.806 13.072 ;
      RECT -20 -20 45.852 13.026 ;
      RECT -20 -20 45.898 12.98 ;
      RECT -20 -20 45.944 12.934 ;
      RECT -20 -20 45.99 12.888 ;
      RECT -20 -20 46.036 12.842 ;
      RECT -20 -20 46.082 12.796 ;
      RECT -20 -20 46.128 12.75 ;
      RECT -20 -20 46.174 12.704 ;
      RECT -20 -20 46.22 12.658 ;
      RECT -20 -20 46.266 12.612 ;
      RECT -20 -20 46.312 12.566 ;
      RECT -20 -20 46.358 12.52 ;
      RECT -20 -20 46.404 12.474 ;
      RECT -20 -20 46.45 12.428 ;
      RECT -20 -20 46.496 12.382 ;
      RECT -20 -20 46.542 12.336 ;
      RECT -20 -20 46.588 12.29 ;
      RECT -20 -20 46.634 12.244 ;
      RECT -20 -20 46.68 12.198 ;
      RECT -20 -20 46.726 12.152 ;
      RECT -20 -20 46.772 12.106 ;
      RECT -20 -20 46.818 12.06 ;
      RECT -20 -20 46.864 12.014 ;
      RECT -20 -20 46.91 11.968 ;
      RECT -20 -20 46.956 11.922 ;
      RECT -20 -20 47.002 11.876 ;
      RECT -20 -20 47.048 11.83 ;
      RECT -20 -20 47.094 11.784 ;
      RECT -20 -20 47.14 11.738 ;
      RECT -20 -20 47.186 11.692 ;
      RECT -20 -20 47.232 11.646 ;
      RECT -20 -20 47.278 11.6 ;
      RECT -20 -20 47.324 11.554 ;
      RECT -20 -20 47.37 11.508 ;
      RECT -20 -20 47.416 11.462 ;
      RECT -20 -20 47.462 11.416 ;
      RECT -20 -20 47.508 11.37 ;
      RECT -20 -20 47.554 11.324 ;
      RECT -20 -20 47.6 11.278 ;
      RECT -20 -20 47.646 11.232 ;
      RECT -20 -20 47.692 11.186 ;
      RECT -20 -20 47.738 11.14 ;
      RECT -20 -20 47.784 11.094 ;
      RECT -20 -20 47.83 11.048 ;
      RECT -20 -20 47.876 11.002 ;
      RECT -20 -20 47.922 10.956 ;
      RECT -20 -20 47.968 10.91 ;
      RECT -20 -20 48.014 10.864 ;
      RECT -20 -20 48.06 10.818 ;
      RECT -20 -20 48.106 10.772 ;
      RECT -20 -20 48.152 10.726 ;
      RECT -20 -20 48.198 10.68 ;
      RECT -20 -20 48.244 10.634 ;
      RECT -20 -20 48.29 10.588 ;
      RECT -20 -20 48.336 10.542 ;
      RECT -20 -20 48.382 10.496 ;
      RECT -20 -20 48.428 10.45 ;
      RECT -20 -20 48.474 10.404 ;
      RECT -20 -20 48.52 10.358 ;
      RECT -20 -20 48.566 10.312 ;
      RECT -20 -20 48.612 10.266 ;
      RECT -20 -20 48.658 10.22 ;
      RECT -20 -20 48.704 10.174 ;
      RECT -20 -20 48.75 10.128 ;
      RECT -20 -20 48.796 10.082 ;
      RECT -20 -20 48.842 10.036 ;
      RECT -20 -20 48.888 9.99 ;
      RECT -20 -20 48.934 9.944 ;
      RECT -20 -20 48.98 9.898 ;
      RECT -20 -20 49.026 9.852 ;
      RECT -20 -20 49.072 9.806 ;
      RECT -20 -20 49.118 9.76 ;
      RECT -20 -20 49.164 9.714 ;
      RECT -20 -20 49.21 9.668 ;
      RECT -20 -20 49.256 9.622 ;
      RECT -20 -20 49.302 9.576 ;
      RECT -20 -20 49.348 9.53 ;
      RECT -20 -20 49.394 9.484 ;
      RECT -20 -20 49.44 9.438 ;
      RECT -20 -20 49.486 9.392 ;
      RECT -20 -20 49.532 9.346 ;
      RECT -20 -20 49.578 9.3 ;
      RECT -20 -20 49.624 9.254 ;
      RECT -20 -20 49.67 9.208 ;
      RECT -20 -20 49.716 9.162 ;
      RECT -20 -20 49.762 9.116 ;
      RECT -20 -20 49.808 9.07 ;
      RECT -20 -20 49.854 9.024 ;
      RECT -20 -20 49.9 8.978 ;
      RECT -20 -20 49.946 8.932 ;
      RECT -20 -20 49.992 8.886 ;
      RECT -20 -20 50.038 8.84 ;
      RECT -20 -20 50.084 8.794 ;
      RECT -20 -20 50.13 8.748 ;
      RECT -20 -20 50.176 8.702 ;
      RECT -20 -20 50.222 8.656 ;
      RECT -20 -20 50.268 8.61 ;
      RECT -20 -20 50.314 8.564 ;
      RECT -20 -20 50.36 8.518 ;
      RECT -20 -20 50.406 8.472 ;
      RECT -20 -20 50.452 8.426 ;
      RECT -20 -20 50.498 8.38 ;
      RECT -20 -20 50.544 8.334 ;
      RECT -20 -20 50.59 8.288 ;
      RECT -20 -20 50.636 8.242 ;
      RECT -20 -20 50.682 8.196 ;
      RECT -20 -20 50.728 8.15 ;
      RECT -20 -20 50.774 8.104 ;
      RECT -20 -20 50.82 8.058 ;
      RECT -20 -20 50.866 8.012 ;
      RECT -20 -20 50.912 7.966 ;
      RECT -20 -20 50.958 7.92 ;
      RECT -20 -20 51.004 7.874 ;
      RECT -20 -20 51.05 7.828 ;
      RECT -20 -20 51.096 7.782 ;
      RECT -20 -20 51.142 7.736 ;
      RECT -20 -20 51.188 7.69 ;
      RECT -20 -20 51.234 7.644 ;
      RECT -20 -20 51.28 7.598 ;
      RECT -20 -20 51.326 7.552 ;
      RECT -20 -20 51.372 7.506 ;
      RECT -20 -20 51.418 7.46 ;
      RECT -20 -20 51.464 7.414 ;
      RECT -20 -20 51.51 7.368 ;
      RECT -20 -20 51.556 7.322 ;
      RECT -20 -20 51.602 7.276 ;
      RECT -20 -20 51.648 7.23 ;
      RECT -20 -20 51.694 7.184 ;
      RECT -20 -20 51.74 7.138 ;
      RECT -20 -20 51.786 7.092 ;
      RECT -20 -20 51.832 7.046 ;
      RECT -20 -20 51.878 7 ;
      RECT -20 -20 51.924 6.954 ;
      RECT -20 -20 51.97 6.908 ;
      RECT -20 -20 52.016 6.862 ;
      RECT -20 -20 52.062 6.816 ;
      RECT -20 -20 52.108 6.77 ;
      RECT -20 -20 52.154 6.724 ;
      RECT -20 -20 52.2 6.678 ;
      RECT -20 -20 52.246 6.632 ;
      RECT -20 -20 52.292 6.586 ;
      RECT -20 -20 52.338 6.54 ;
      RECT -20 -20 52.384 6.494 ;
      RECT -20 -20 52.43 6.448 ;
      RECT -20 -20 52.476 6.402 ;
      RECT -20 -20 52.522 6.356 ;
      RECT -20 -20 52.568 6.31 ;
      RECT -20 -20 52.614 6.264 ;
      RECT -20 -20 52.66 6.218 ;
      RECT -20 -20 52.706 6.172 ;
      RECT -20 -20 52.752 6.126 ;
      RECT -20 -20 52.798 6.08 ;
      RECT -20 -20 52.844 6.034 ;
      RECT -20 -20 52.89 5.988 ;
      RECT -20 -20 52.936 5.942 ;
      RECT -20 -20 52.982 5.896 ;
      RECT -20 -20 53.028 5.85 ;
      RECT -20 -20 53.074 5.804 ;
      RECT -20 -20 53.12 5.758 ;
      RECT -20 -20 53.166 5.712 ;
      RECT -20 -20 53.212 5.666 ;
      RECT -20 -20 53.258 5.62 ;
      RECT -20 -20 53.304 5.574 ;
      RECT -20 -20 53.35 5.528 ;
      RECT -20 -20 53.396 5.482 ;
      RECT -20 -20 53.442 5.436 ;
      RECT -20 -20 53.488 5.39 ;
      RECT -20 -20 53.534 5.344 ;
      RECT -20 -20 53.58 5.298 ;
      RECT -20 -20 53.626 5.252 ;
      RECT -20 -20 53.672 5.206 ;
      RECT -20 -20 53.718 5.16 ;
      RECT -20 -20 53.764 5.114 ;
      RECT -20 -20 53.81 5.068 ;
      RECT -20 -20 53.856 5.022 ;
      RECT -20 -20 53.902 4.976 ;
      RECT -20 -20 53.948 4.93 ;
      RECT -20 -20 53.994 4.884 ;
      RECT -20 -20 54.04 4.838 ;
      RECT -20 -20 54.086 4.792 ;
      RECT -20 -20 54.132 4.746 ;
      RECT -20 -20 54.178 4.7 ;
      RECT -20 -20 54.224 4.654 ;
      RECT -20 -20 54.27 4.608 ;
      RECT -20 -20 54.316 4.562 ;
      RECT -20 -20 54.362 4.516 ;
      RECT -20 -20 54.408 4.47 ;
      RECT -20 -20 54.454 4.424 ;
      RECT -20 -20 54.5 4.378 ;
      RECT -20 -20 54.546 4.332 ;
      RECT -20 -20 54.592 4.286 ;
      RECT -20 -20 54.638 4.24 ;
      RECT -20 -20 54.684 4.194 ;
      RECT -20 -20 54.73 4.148 ;
      RECT -20 -20 54.776 4.102 ;
      RECT -20 -20 54.822 4.056 ;
      RECT -20 -20 54.868 4.01 ;
      RECT -20 -20 54.914 3.964 ;
      RECT -20 -20 54.96 3.918 ;
      RECT -20 -20 55.006 3.872 ;
      RECT -20 -20 55.052 3.826 ;
      RECT -20 -20 55.098 3.78 ;
      RECT -20 -20 55.144 3.734 ;
      RECT -20 -20 55.19 3.688 ;
      RECT -20 -20 55.236 3.642 ;
      RECT -20 -20 55.282 3.596 ;
      RECT -20 -20 55.328 3.55 ;
      RECT -20 -20 55.374 3.504 ;
      RECT -20 -20 55.42 3.458 ;
      RECT -20 -20 55.466 3.412 ;
      RECT -20 -20 55.512 3.366 ;
      RECT -20 -20 55.558 3.32 ;
      RECT -20 -20 55.604 3.274 ;
      RECT -20 -20 55.65 3.228 ;
      RECT -20 -20 55.685 3.187 ;
      RECT -20 -20 110 3.17 ;
      RECT 15.83 61.287 16.67 110 ;
      RECT 15.83 61.287 16.716 62.412 ;
      RECT 15.83 61.287 16.762 62.366 ;
      RECT 15.83 61.287 16.808 62.32 ;
      RECT 15.83 61.287 16.854 62.274 ;
      RECT 15.83 61.287 16.9 62.228 ;
      RECT 15.83 61.287 16.946 62.182 ;
      RECT 15.83 61.287 16.992 62.136 ;
      RECT 15.83 61.287 17.038 62.09 ;
      RECT 15.83 61.287 17.084 62.044 ;
      RECT 15.83 61.287 17.13 61.998 ;
      RECT 15.83 61.287 17.176 61.952 ;
      RECT 15.83 61.287 17.222 61.906 ;
      RECT 15.83 61.287 17.268 61.86 ;
      RECT 15.83 61.287 17.314 61.814 ;
      RECT 15.83 61.287 17.36 61.768 ;
      RECT 15.83 61.287 17.406 61.722 ;
      RECT 15.83 61.287 17.452 61.676 ;
      RECT 15.83 61.287 17.498 61.63 ;
      RECT 15.83 61.287 17.544 61.584 ;
      RECT 15.83 61.287 17.59 61.538 ;
      RECT 15.83 61.287 17.636 61.492 ;
      RECT 15.83 61.287 17.682 61.446 ;
      RECT 15.83 61.287 17.728 61.4 ;
      RECT 15.83 61.287 17.774 61.354 ;
      RECT 15.876 61.241 17.82 61.308 ;
      RECT 17.762 59.355 17.82 61.308 ;
      RECT 15.922 61.195 17.866 61.262 ;
      RECT 17.808 59.309 17.866 61.262 ;
      RECT 15.968 61.149 17.912 61.216 ;
      RECT 17.854 59.263 17.912 61.216 ;
      RECT 16.014 61.103 17.958 61.17 ;
      RECT 17.9 59.217 17.958 61.17 ;
      RECT 16.06 61.057 18.004 61.124 ;
      RECT 17.946 59.171 18.004 61.124 ;
      RECT 16.106 61.011 18.05 61.078 ;
      RECT 17.992 59.125 18.05 61.078 ;
      RECT 16.152 60.965 18.096 61.032 ;
      RECT 18.038 59.079 18.096 61.032 ;
      RECT 16.198 60.919 18.142 60.986 ;
      RECT 18.084 59.033 18.142 60.986 ;
      RECT 16.244 60.873 18.188 60.94 ;
      RECT 18.13 58.987 18.188 60.94 ;
      RECT 16.29 60.827 18.234 60.894 ;
      RECT 18.176 58.941 18.234 60.894 ;
      RECT 16.336 60.781 18.28 60.848 ;
      RECT 18.222 58.895 18.28 60.848 ;
      RECT 16.382 60.735 18.326 60.802 ;
      RECT 18.268 58.849 18.326 60.802 ;
      RECT 16.428 60.689 18.372 60.756 ;
      RECT 18.314 58.803 18.372 60.756 ;
      RECT 16.474 60.643 18.418 60.71 ;
      RECT 18.36 58.757 18.418 60.71 ;
      RECT 16.52 60.597 18.464 60.664 ;
      RECT 18.406 58.711 18.464 60.664 ;
      RECT 16.566 60.551 18.51 60.618 ;
      RECT 18.452 58.665 18.51 60.618 ;
      RECT 16.612 60.505 18.556 60.572 ;
      RECT 18.498 58.619 18.556 60.572 ;
      RECT 16.658 60.459 18.602 60.526 ;
      RECT 18.544 58.573 18.602 60.526 ;
      RECT 16.704 60.413 18.648 60.48 ;
      RECT 18.59 58.527 18.648 60.48 ;
      RECT 16.75 60.367 18.694 60.434 ;
      RECT 18.636 58.481 18.694 60.434 ;
      RECT 16.796 60.321 18.74 60.388 ;
      RECT 18.682 58.435 18.74 60.388 ;
      RECT 16.842 60.275 18.786 60.342 ;
      RECT 18.728 58.389 18.786 60.342 ;
      RECT 16.888 60.229 18.832 60.296 ;
      RECT 18.774 58.343 18.832 60.296 ;
      RECT 16.934 60.183 18.878 60.25 ;
      RECT 18.82 58.297 18.878 60.25 ;
      RECT 16.98 60.137 18.924 60.204 ;
      RECT 18.866 58.251 18.924 60.204 ;
      RECT 17.026 60.091 18.97 60.158 ;
      RECT 18.912 58.205 18.97 60.158 ;
      RECT 17.072 60.045 19.016 60.112 ;
      RECT 18.958 58.159 19.016 60.112 ;
      RECT 17.118 59.999 19.062 60.066 ;
      RECT 19.004 58.113 19.062 60.066 ;
      RECT 17.164 59.953 19.108 60.02 ;
      RECT 19.05 58.067 19.108 60.02 ;
      RECT 17.21 59.907 19.154 59.974 ;
      RECT 19.096 58.021 19.154 59.974 ;
      RECT 17.256 59.861 19.2 59.928 ;
      RECT 19.142 57.975 19.2 59.928 ;
      RECT 17.302 59.815 19.246 59.882 ;
      RECT 19.188 57.929 19.246 59.882 ;
      RECT 17.348 59.769 19.292 59.836 ;
      RECT 19.234 57.883 19.292 59.836 ;
      RECT 17.394 59.723 19.338 59.79 ;
      RECT 19.28 57.837 19.338 59.79 ;
      RECT 17.44 59.677 19.384 59.744 ;
      RECT 19.326 57.791 19.384 59.744 ;
      RECT 17.486 59.631 19.43 59.698 ;
      RECT 19.372 57.745 19.43 59.698 ;
      RECT 17.532 59.585 19.476 59.652 ;
      RECT 19.418 57.699 19.476 59.652 ;
      RECT 17.578 59.539 19.522 59.606 ;
      RECT 19.464 57.653 19.522 59.606 ;
      RECT 17.624 59.493 19.568 59.56 ;
      RECT 19.51 57.607 19.568 59.56 ;
      RECT 17.67 59.447 19.614 59.514 ;
      RECT 19.556 57.561 19.614 59.514 ;
      RECT 17.716 59.401 19.66 59.468 ;
      RECT 19.602 57.515 19.66 59.468 ;
      RECT 19.648 57.469 19.706 59.422 ;
      RECT 19.694 57.423 19.752 59.376 ;
      RECT 19.74 57.377 19.798 59.33 ;
      RECT 19.786 57.331 19.844 59.284 ;
      RECT 19.832 57.285 19.89 59.238 ;
      RECT 19.878 57.239 19.936 59.192 ;
      RECT 19.924 57.193 19.982 59.146 ;
      RECT 19.97 57.147 20.028 59.1 ;
      RECT 20.016 57.101 20.074 59.054 ;
      RECT 20.062 57.055 20.12 59.008 ;
      RECT 20.108 57.009 20.166 58.962 ;
      RECT 20.154 56.963 20.212 58.916 ;
      RECT 20.2 56.917 20.258 58.87 ;
      RECT 20.246 56.871 20.304 58.824 ;
      RECT 20.292 56.825 20.35 58.778 ;
      RECT 20.338 56.779 20.396 58.732 ;
      RECT 20.384 56.733 20.442 58.686 ;
      RECT 20.43 56.687 20.488 58.64 ;
      RECT 20.476 56.641 20.534 58.594 ;
      RECT 20.522 56.595 20.58 58.548 ;
      RECT 20.568 56.549 20.626 58.502 ;
      RECT 20.614 56.503 20.672 58.456 ;
      RECT 20.66 56.457 20.718 58.41 ;
      RECT 20.706 56.411 20.764 58.364 ;
      RECT 20.752 56.365 20.81 58.318 ;
      RECT 20.798 56.319 20.856 58.272 ;
      RECT 20.844 56.273 20.902 58.226 ;
      RECT 20.89 56.227 20.948 58.18 ;
      RECT 20.936 56.181 20.994 58.134 ;
      RECT 20.982 56.135 21.04 58.088 ;
      RECT 21.028 56.089 21.086 58.042 ;
      RECT 21.074 56.043 21.132 57.996 ;
      RECT 21.12 55.997 21.178 57.95 ;
      RECT 21.166 55.951 21.224 57.904 ;
      RECT 21.212 55.905 21.27 57.858 ;
      RECT 21.258 55.859 21.316 57.812 ;
      RECT 21.304 55.813 21.362 57.766 ;
      RECT 21.35 55.767 21.408 57.72 ;
      RECT 21.396 55.721 21.454 57.674 ;
      RECT 21.442 55.675 21.5 57.628 ;
      RECT 21.488 55.629 21.546 57.582 ;
      RECT 21.534 55.583 21.592 57.536 ;
      RECT 21.58 55.537 21.638 57.49 ;
      RECT 21.626 55.491 21.684 57.444 ;
      RECT 21.672 55.445 21.73 57.398 ;
      RECT 21.718 55.399 21.776 57.352 ;
      RECT 21.764 55.353 21.822 57.306 ;
      RECT 21.81 55.307 21.868 57.26 ;
      RECT 21.856 55.261 21.914 57.214 ;
      RECT 21.902 55.215 21.96 57.168 ;
      RECT 21.948 55.169 22.006 57.122 ;
      RECT 21.994 55.123 22.052 57.076 ;
      RECT 22.04 55.077 22.098 57.03 ;
      RECT 22.086 55.031 22.144 56.984 ;
      RECT 22.132 54.985 22.19 56.938 ;
      RECT 22.178 54.939 22.236 56.892 ;
      RECT 22.224 54.893 22.282 56.846 ;
      RECT 22.27 54.847 22.328 56.8 ;
      RECT 22.316 54.801 22.374 56.754 ;
      RECT 22.362 54.755 22.42 56.708 ;
      RECT 22.408 54.709 22.466 56.662 ;
      RECT 22.454 54.663 22.512 56.616 ;
      RECT 22.5 54.617 22.558 56.57 ;
      RECT 22.546 54.571 22.604 56.524 ;
      RECT 22.592 54.525 22.65 56.478 ;
      RECT 22.638 54.479 22.696 56.432 ;
      RECT 22.684 54.433 22.742 56.386 ;
      RECT 22.73 54.387 22.788 56.34 ;
      RECT 22.776 54.341 22.834 56.294 ;
      RECT 22.822 54.295 22.88 56.248 ;
      RECT 22.868 54.249 22.926 56.202 ;
      RECT 22.914 54.203 22.972 56.156 ;
      RECT 22.96 54.157 23.018 56.11 ;
      RECT 23.006 54.111 23.064 56.064 ;
      RECT 23.052 54.065 23.11 56.018 ;
      RECT 23.098 54.019 23.156 55.972 ;
      RECT 23.144 53.973 23.202 55.926 ;
      RECT 23.19 53.927 23.248 55.88 ;
      RECT 23.236 53.881 23.294 55.834 ;
      RECT 23.282 53.835 23.34 55.788 ;
      RECT 23.328 53.789 23.386 55.742 ;
      RECT 23.374 53.743 23.432 55.696 ;
      RECT 23.42 53.697 23.478 55.65 ;
      RECT 23.466 53.651 23.524 55.604 ;
      RECT 23.512 53.605 23.57 55.558 ;
      RECT 23.558 53.559 23.616 55.512 ;
      RECT 23.604 53.513 23.662 55.466 ;
      RECT 23.65 53.467 23.708 55.42 ;
      RECT 23.696 53.421 23.754 55.374 ;
      RECT 23.742 53.375 23.8 55.328 ;
      RECT 23.788 53.329 23.846 55.282 ;
      RECT 23.834 53.283 23.892 55.236 ;
      RECT 23.88 53.237 23.938 55.19 ;
      RECT 23.926 53.191 23.984 55.144 ;
      RECT 23.972 53.145 24.03 55.098 ;
      RECT 24.018 53.099 24.076 55.052 ;
      RECT 24.064 53.053 24.122 55.006 ;
      RECT 24.11 53.007 24.168 54.96 ;
      RECT 24.156 52.961 24.214 54.914 ;
      RECT 24.202 52.915 24.26 54.868 ;
      RECT 24.248 52.869 24.306 54.822 ;
      RECT 24.294 52.823 24.352 54.776 ;
      RECT 24.34 52.777 24.398 54.73 ;
      RECT 24.386 52.731 24.444 54.684 ;
      RECT 24.432 52.685 24.49 54.638 ;
      RECT 24.478 52.639 24.536 54.592 ;
      RECT 24.524 52.593 24.582 54.546 ;
      RECT 24.57 52.547 24.628 54.5 ;
      RECT 24.616 52.501 24.674 54.454 ;
      RECT 24.662 52.455 24.72 54.408 ;
      RECT 24.708 52.409 24.766 54.362 ;
      RECT 24.754 52.363 24.812 54.316 ;
      RECT 24.8 52.317 24.858 54.27 ;
      RECT 24.846 52.271 24.904 54.224 ;
      RECT 24.892 52.225 24.95 54.178 ;
      RECT 24.938 52.179 24.996 54.132 ;
      RECT 24.984 52.133 25.042 54.086 ;
      RECT 25.03 52.087 25.088 54.04 ;
      RECT 25.076 52.041 25.134 53.994 ;
      RECT 25.122 51.995 25.18 53.948 ;
      RECT 25.168 51.949 25.226 53.902 ;
      RECT 25.214 51.903 25.272 53.856 ;
      RECT 25.26 51.857 25.318 53.81 ;
      RECT 25.306 51.811 25.364 53.764 ;
      RECT 25.352 51.765 25.41 53.718 ;
      RECT 25.398 51.719 25.456 53.672 ;
      RECT 25.444 51.673 25.502 53.626 ;
      RECT 25.49 51.627 25.548 53.58 ;
      RECT 25.536 51.581 25.594 53.534 ;
      RECT 25.582 51.535 25.64 53.488 ;
      RECT 25.628 51.489 25.686 53.442 ;
      RECT 25.674 51.443 25.732 53.396 ;
      RECT 25.72 51.397 25.778 53.35 ;
      RECT 25.766 51.351 25.824 53.304 ;
      RECT 25.812 51.305 25.87 53.258 ;
      RECT 25.858 51.259 25.916 53.212 ;
      RECT 25.904 51.213 25.962 53.166 ;
      RECT 25.95 51.167 26.008 53.12 ;
      RECT 25.996 51.121 26.054 53.074 ;
      RECT 26.042 51.075 26.1 53.028 ;
      RECT 26.088 51.029 26.146 52.982 ;
      RECT 26.134 50.983 26.192 52.936 ;
      RECT 26.18 50.937 26.238 52.89 ;
      RECT 26.226 50.891 26.284 52.844 ;
      RECT 26.272 50.845 26.33 52.798 ;
      RECT 26.318 50.799 26.376 52.752 ;
      RECT 26.364 50.753 26.422 52.706 ;
      RECT 26.41 50.707 26.468 52.66 ;
      RECT 26.456 50.661 26.514 52.614 ;
      RECT 26.502 50.615 26.56 52.568 ;
      RECT 26.548 50.569 26.606 52.522 ;
      RECT 26.594 50.523 26.652 52.476 ;
      RECT 26.64 50.477 26.698 52.43 ;
      RECT 26.686 50.431 26.744 52.384 ;
      RECT 26.732 50.385 26.79 52.338 ;
      RECT 26.778 50.339 26.836 52.292 ;
      RECT 26.824 50.293 26.882 52.246 ;
      RECT 26.87 50.247 26.928 52.2 ;
      RECT 26.916 50.201 26.974 52.154 ;
      RECT 26.962 50.155 27.02 52.108 ;
      RECT 27.008 50.109 27.066 52.062 ;
      RECT 27.054 50.063 27.112 52.016 ;
      RECT 27.1 50.017 27.158 51.97 ;
      RECT 27.146 49.971 27.204 51.924 ;
      RECT 27.192 49.925 27.25 51.878 ;
      RECT 27.238 49.879 27.296 51.832 ;
      RECT 27.284 49.833 27.342 51.786 ;
      RECT 27.33 49.787 27.388 51.74 ;
      RECT 27.376 49.741 27.434 51.694 ;
      RECT 27.422 49.695 27.48 51.648 ;
      RECT 27.468 49.649 27.526 51.602 ;
      RECT 27.514 49.603 27.572 51.556 ;
      RECT 27.56 49.557 27.618 51.51 ;
      RECT 27.606 49.511 27.664 51.464 ;
      RECT 27.652 49.465 27.71 51.418 ;
      RECT 27.698 49.419 27.756 51.372 ;
      RECT 27.744 49.373 27.802 51.326 ;
      RECT 27.79 49.327 27.848 51.28 ;
      RECT 27.836 49.281 27.894 51.234 ;
      RECT 27.882 49.235 27.94 51.188 ;
      RECT 27.928 49.189 27.986 51.142 ;
      RECT 27.974 49.143 28.032 51.096 ;
      RECT 28.02 49.097 28.078 51.05 ;
      RECT 28.066 49.051 28.124 51.004 ;
      RECT 28.112 49.005 28.17 50.958 ;
      RECT 28.158 48.959 28.216 50.912 ;
      RECT 28.204 48.913 28.262 50.866 ;
      RECT 28.25 48.867 28.308 50.82 ;
      RECT 28.296 48.821 28.354 50.774 ;
      RECT 28.342 48.775 28.4 50.728 ;
      RECT 28.388 48.729 28.446 50.682 ;
      RECT 28.434 48.683 28.492 50.636 ;
      RECT 28.48 48.637 28.538 50.59 ;
      RECT 28.526 48.591 28.584 50.544 ;
      RECT 28.572 48.545 28.63 50.498 ;
      RECT 28.618 48.499 28.67 50.455 ;
      RECT 28.664 48.453 28.716 50.412 ;
      RECT 28.71 48.407 28.762 50.366 ;
      RECT 28.756 48.361 28.808 50.32 ;
      RECT 28.802 48.315 28.854 50.274 ;
      RECT 28.848 48.269 28.9 50.228 ;
      RECT 28.894 48.223 28.946 50.182 ;
      RECT 28.94 48.177 28.992 50.136 ;
      RECT 28.986 48.131 29.038 50.09 ;
      RECT 29.032 48.085 29.084 50.044 ;
      RECT 29.078 48.039 29.13 49.998 ;
      RECT 29.124 47.993 29.176 49.952 ;
      RECT 29.17 47.947 29.222 49.906 ;
      RECT 29.216 47.901 29.268 49.86 ;
      RECT 29.262 47.855 29.314 49.814 ;
      RECT 29.308 47.809 29.36 49.768 ;
      RECT 29.354 47.763 29.406 49.722 ;
      RECT 29.4 47.717 29.452 49.676 ;
      RECT 29.446 47.671 29.498 49.63 ;
      RECT 29.492 47.625 29.544 49.584 ;
      RECT 29.538 47.579 29.59 49.538 ;
      RECT 29.584 47.533 29.636 49.492 ;
      RECT 29.63 47.487 29.682 49.446 ;
      RECT 29.676 47.441 29.728 49.4 ;
      RECT 29.722 47.395 29.774 49.354 ;
      RECT 29.768 47.349 29.82 49.308 ;
      RECT 29.814 47.303 29.866 49.262 ;
      RECT 29.86 47.257 29.912 49.216 ;
      RECT 29.906 47.211 29.958 49.17 ;
      RECT 29.952 47.165 30.004 49.124 ;
      RECT 29.998 47.119 30.05 49.078 ;
      RECT 30.044 47.073 30.096 49.032 ;
      RECT 30.09 47.027 30.142 48.986 ;
      RECT 30.136 46.981 30.188 48.94 ;
      RECT 30.182 46.935 30.234 48.894 ;
      RECT 30.228 46.889 30.28 48.848 ;
      RECT 30.274 46.843 30.326 48.802 ;
      RECT 30.32 46.797 30.372 48.756 ;
      RECT 30.366 46.751 30.418 48.71 ;
      RECT 30.412 46.705 30.464 48.664 ;
      RECT 30.458 46.659 30.51 48.618 ;
      RECT 30.504 46.613 30.556 48.572 ;
      RECT 30.55 46.567 30.602 48.526 ;
      RECT 30.596 46.521 30.648 48.48 ;
      RECT 30.642 46.475 30.694 48.434 ;
      RECT 30.688 46.429 30.74 48.388 ;
      RECT 30.734 46.383 30.786 48.342 ;
      RECT 30.78 46.337 30.832 48.296 ;
      RECT 30.826 46.291 30.878 48.25 ;
      RECT 30.872 46.245 30.924 48.204 ;
      RECT 30.918 46.199 30.97 48.158 ;
      RECT 30.964 46.153 31.016 48.112 ;
      RECT 31.01 46.107 31.062 48.066 ;
      RECT 31.056 46.061 31.108 48.02 ;
      RECT 31.102 46.015 31.154 47.974 ;
      RECT 31.148 45.969 31.2 47.928 ;
      RECT 31.194 45.923 31.246 47.882 ;
      RECT 31.24 45.877 31.292 47.836 ;
      RECT 31.286 45.831 31.338 47.79 ;
      RECT 31.332 45.785 31.384 47.744 ;
      RECT 31.378 45.739 31.43 47.698 ;
      RECT 31.424 45.693 31.476 47.652 ;
      RECT 31.47 45.647 31.522 47.606 ;
      RECT 31.516 45.601 31.568 47.56 ;
      RECT 31.562 45.555 31.614 47.514 ;
      RECT 31.608 45.509 31.66 47.468 ;
      RECT 31.654 45.463 31.706 47.422 ;
      RECT 31.7 45.417 31.752 47.376 ;
      RECT 31.746 45.371 31.798 47.33 ;
      RECT 31.792 45.325 31.844 47.284 ;
      RECT 31.838 45.279 31.89 47.238 ;
      RECT 31.884 45.233 31.936 47.192 ;
      RECT 31.93 45.187 31.982 47.146 ;
      RECT 31.976 45.141 32.028 47.1 ;
      RECT 32.022 45.095 32.074 47.054 ;
      RECT 32.068 45.049 32.12 47.008 ;
      RECT 32.114 45.003 32.166 46.962 ;
      RECT 32.16 44.957 32.212 46.916 ;
      RECT 32.206 44.911 32.258 46.87 ;
      RECT 32.252 44.865 32.304 46.824 ;
      RECT 32.298 44.819 32.35 46.778 ;
      RECT 32.344 44.773 32.396 46.732 ;
      RECT 32.39 44.727 32.442 46.686 ;
      RECT 32.436 44.681 32.488 46.64 ;
      RECT 32.482 44.635 32.534 46.594 ;
      RECT 32.528 44.589 32.58 46.548 ;
      RECT 32.574 44.543 32.626 46.502 ;
      RECT 32.62 44.497 32.672 46.456 ;
      RECT 32.666 44.451 32.718 46.41 ;
      RECT 32.712 44.405 32.764 46.364 ;
      RECT 32.758 44.359 32.81 46.318 ;
      RECT 32.804 44.313 32.856 46.272 ;
      RECT 32.85 44.267 32.902 46.226 ;
      RECT 32.896 44.221 32.948 46.18 ;
      RECT 32.942 44.175 32.994 46.134 ;
      RECT 32.988 44.129 33.04 46.088 ;
      RECT 33.034 44.083 33.086 46.042 ;
      RECT 33.08 44.037 33.132 45.996 ;
      RECT 33.126 43.991 33.178 45.95 ;
      RECT 33.172 43.945 33.224 45.904 ;
      RECT 33.218 43.899 33.27 45.858 ;
      RECT 33.264 43.853 33.316 45.812 ;
      RECT 33.31 43.807 33.362 45.766 ;
      RECT 33.356 43.761 33.408 45.72 ;
      RECT 33.402 43.715 33.454 45.674 ;
      RECT 33.448 43.669 33.5 45.628 ;
      RECT 33.494 43.623 33.546 45.582 ;
      RECT 33.54 43.577 33.592 45.536 ;
      RECT 33.586 43.531 33.638 45.49 ;
      RECT 33.632 43.485 33.684 45.444 ;
      RECT 33.678 43.439 33.73 45.398 ;
      RECT 33.724 43.393 33.776 45.352 ;
      RECT 33.77 43.347 33.822 45.306 ;
      RECT 33.816 43.301 33.868 45.26 ;
      RECT 33.862 43.255 33.914 45.214 ;
      RECT 33.908 43.209 33.96 45.168 ;
      RECT 33.954 43.163 34.006 45.122 ;
      RECT 34 43.117 34.052 45.076 ;
      RECT 34.046 43.071 34.098 45.03 ;
      RECT 34.092 43.025 34.144 44.984 ;
      RECT 34.138 42.979 34.19 44.938 ;
      RECT 34.184 42.933 34.236 44.892 ;
      RECT 34.23 42.887 34.282 44.846 ;
      RECT 34.276 42.841 34.328 44.8 ;
      RECT 34.322 42.795 34.374 44.754 ;
      RECT 34.368 42.749 34.42 44.708 ;
      RECT 34.414 42.703 34.466 44.662 ;
      RECT 34.46 42.657 34.512 44.616 ;
      RECT 34.506 42.611 34.558 44.57 ;
      RECT 34.552 42.565 34.604 44.524 ;
      RECT 34.598 42.519 34.65 44.478 ;
      RECT 34.644 42.473 34.696 44.432 ;
      RECT 34.69 42.427 34.742 44.386 ;
      RECT 34.736 42.381 34.788 44.34 ;
      RECT 34.782 42.335 34.834 44.294 ;
      RECT 34.828 42.289 34.88 44.248 ;
      RECT 34.874 42.243 34.926 44.202 ;
      RECT 34.92 42.197 34.972 44.156 ;
      RECT 34.966 42.151 35.018 44.11 ;
      RECT 35.012 42.105 35.064 44.064 ;
      RECT 35.058 42.059 35.11 44.018 ;
      RECT 35.104 42.013 35.156 43.972 ;
      RECT 35.15 41.967 35.202 43.926 ;
      RECT 35.196 41.921 35.248 43.88 ;
      RECT 35.242 41.875 35.294 43.834 ;
      RECT 35.288 41.829 35.34 43.788 ;
      RECT 35.334 41.783 35.386 43.742 ;
      RECT 35.38 41.737 35.432 43.696 ;
      RECT 35.426 41.691 35.478 43.65 ;
      RECT 35.472 41.645 35.524 43.604 ;
      RECT 35.518 41.599 35.57 43.558 ;
      RECT 35.564 41.553 35.616 43.512 ;
      RECT 35.61 41.507 35.662 43.466 ;
      RECT 35.656 41.461 35.708 43.42 ;
      RECT 35.702 41.415 35.754 43.374 ;
      RECT 35.748 41.369 35.8 43.328 ;
      RECT 35.794 41.323 35.846 43.282 ;
      RECT 35.84 41.277 35.892 43.236 ;
      RECT 35.886 41.231 35.938 43.19 ;
      RECT 35.932 41.185 35.984 43.144 ;
      RECT 35.978 41.139 36.03 43.098 ;
      RECT 36.024 41.093 36.076 43.052 ;
      RECT 36.07 41.047 36.122 43.006 ;
      RECT 36.116 41.001 36.168 42.96 ;
      RECT 36.162 40.955 36.214 42.914 ;
      RECT 36.208 40.909 36.26 42.868 ;
      RECT 36.254 40.863 36.306 42.822 ;
      RECT 36.3 40.817 36.352 42.776 ;
      RECT 36.346 40.771 36.398 42.73 ;
      RECT 36.392 40.725 36.444 42.684 ;
      RECT 36.438 40.679 36.49 42.638 ;
      RECT 36.484 40.633 36.536 42.592 ;
      RECT 36.53 40.587 36.582 42.546 ;
      RECT 36.576 40.541 36.628 42.5 ;
      RECT 36.622 40.495 36.674 42.454 ;
      RECT 36.668 40.449 36.72 42.408 ;
      RECT 36.714 40.403 36.766 42.362 ;
      RECT 36.76 40.357 36.812 42.316 ;
      RECT 36.806 40.311 36.858 42.27 ;
      RECT 36.852 40.265 36.904 42.224 ;
      RECT 36.898 40.219 36.95 42.178 ;
      RECT 36.944 40.173 36.996 42.132 ;
      RECT 36.99 40.127 37.042 42.086 ;
      RECT 37.036 40.081 37.088 42.04 ;
      RECT 37.082 40.035 37.134 41.994 ;
      RECT 37.128 39.989 37.18 41.948 ;
      RECT 37.174 39.943 37.226 41.902 ;
      RECT 37.22 39.897 37.272 41.856 ;
      RECT 37.266 39.851 37.318 41.81 ;
      RECT 37.312 39.805 37.364 41.764 ;
      RECT 37.358 39.759 37.41 41.718 ;
      RECT 37.404 39.713 37.456 41.672 ;
      RECT 37.45 39.667 37.502 41.626 ;
      RECT 37.496 39.621 37.548 41.58 ;
      RECT 37.542 39.575 37.594 41.534 ;
      RECT 37.588 39.529 37.64 41.488 ;
      RECT 37.634 39.483 37.686 41.442 ;
      RECT 37.68 39.437 37.732 41.396 ;
      RECT 37.726 39.391 37.778 41.35 ;
      RECT 37.772 39.345 37.824 41.304 ;
      RECT 37.818 39.299 37.87 41.258 ;
      RECT 37.864 39.253 37.916 41.212 ;
      RECT 37.91 39.207 37.962 41.166 ;
      RECT 37.956 39.161 38.008 41.12 ;
      RECT 38.002 39.115 38.054 41.074 ;
      RECT 38.048 39.069 38.1 41.028 ;
      RECT 38.094 39.023 38.146 40.982 ;
      RECT 38.14 38.977 38.192 40.936 ;
      RECT 38.186 38.931 38.238 40.89 ;
      RECT 38.232 38.885 38.284 40.844 ;
      RECT 38.278 38.839 38.33 40.798 ;
      RECT 38.324 38.793 38.376 40.752 ;
      RECT 38.37 38.747 38.422 40.706 ;
      RECT 38.416 38.701 38.468 40.66 ;
      RECT 38.462 38.655 38.514 40.614 ;
      RECT 38.508 38.609 38.56 40.568 ;
      RECT 38.554 38.563 38.606 40.522 ;
      RECT 38.6 38.517 38.652 40.476 ;
      RECT 38.646 38.471 38.698 40.43 ;
      RECT 38.692 38.425 38.744 40.384 ;
      RECT 38.738 38.379 38.79 40.338 ;
      RECT 38.784 38.333 38.836 40.292 ;
      RECT 38.83 38.287 38.882 40.246 ;
      RECT 38.876 38.241 38.928 40.2 ;
      RECT 38.922 38.195 38.974 40.154 ;
      RECT 38.968 38.149 39.02 40.108 ;
      RECT 39.014 38.103 39.066 40.062 ;
      RECT 39.06 38.057 39.112 40.016 ;
      RECT 39.106 38.011 39.158 39.97 ;
      RECT 39.152 37.965 39.204 39.924 ;
      RECT 39.198 37.919 39.25 39.878 ;
      RECT 39.244 37.873 39.296 39.832 ;
      RECT 39.29 37.827 39.342 39.786 ;
      RECT 39.336 37.781 39.388 39.74 ;
      RECT 39.382 37.735 39.434 39.694 ;
      RECT 39.428 37.689 39.48 39.648 ;
      RECT 39.474 37.643 39.526 39.602 ;
      RECT 39.52 37.597 39.572 39.556 ;
      RECT 39.566 37.551 39.618 39.51 ;
      RECT 39.612 37.505 39.664 39.464 ;
      RECT 39.658 37.459 39.71 39.418 ;
      RECT 39.704 37.413 39.756 39.372 ;
      RECT 39.75 37.367 39.802 39.326 ;
      RECT 39.796 37.321 39.848 39.28 ;
      RECT 39.842 37.275 39.894 39.234 ;
      RECT 39.888 37.229 39.94 39.188 ;
      RECT 39.934 37.183 39.986 39.142 ;
      RECT 39.98 37.137 40.032 39.096 ;
      RECT 40.026 37.091 40.078 39.05 ;
      RECT 40.072 37.045 40.124 39.004 ;
      RECT 40.118 36.999 40.17 38.958 ;
      RECT 40.164 36.953 40.216 38.912 ;
      RECT 40.21 36.907 40.262 38.866 ;
      RECT 40.256 36.861 40.308 38.82 ;
      RECT 40.302 36.815 40.354 38.774 ;
      RECT 40.348 36.769 40.4 38.728 ;
      RECT 40.394 36.723 40.446 38.682 ;
      RECT 40.44 36.677 40.492 38.636 ;
      RECT 40.486 36.631 40.538 38.59 ;
      RECT 40.532 36.585 40.584 38.544 ;
      RECT 40.578 36.539 40.63 38.498 ;
      RECT 40.624 36.493 40.676 38.452 ;
      RECT 40.67 36.447 40.722 38.406 ;
      RECT 40.716 36.401 40.768 38.36 ;
      RECT 40.762 36.355 40.814 38.314 ;
      RECT 40.808 36.309 40.86 38.268 ;
      RECT 40.854 36.263 40.906 38.222 ;
      RECT 40.9 36.217 40.952 38.176 ;
      RECT 40.946 36.171 40.998 38.13 ;
      RECT 40.992 36.125 41.044 38.084 ;
      RECT 41.038 36.079 41.09 38.038 ;
      RECT 41.084 36.033 41.136 37.992 ;
      RECT 41.13 35.987 41.182 37.946 ;
      RECT 41.176 35.941 41.228 37.9 ;
      RECT 41.222 35.895 41.274 37.854 ;
      RECT 41.268 35.849 41.32 37.808 ;
      RECT 41.314 35.803 41.366 37.762 ;
      RECT 41.36 35.757 41.412 37.716 ;
      RECT 41.406 35.711 41.458 37.67 ;
      RECT 41.452 35.665 41.504 37.624 ;
      RECT 41.498 35.619 41.55 37.578 ;
      RECT 41.544 35.573 41.596 37.532 ;
      RECT 41.59 35.527 41.642 37.486 ;
      RECT 41.636 35.481 41.688 37.44 ;
      RECT 41.682 35.435 41.734 37.394 ;
      RECT 41.728 35.389 41.78 37.348 ;
      RECT 41.774 35.343 41.826 37.302 ;
      RECT 41.82 35.297 41.872 37.256 ;
      RECT 41.866 35.251 41.918 37.21 ;
      RECT 41.912 35.205 41.964 37.164 ;
      RECT 41.958 35.159 42.01 37.118 ;
      RECT 42.004 35.113 42.056 37.072 ;
      RECT 42.05 35.067 42.102 37.026 ;
      RECT 42.096 35.021 42.148 36.98 ;
      RECT 42.142 34.975 42.194 36.934 ;
      RECT 42.188 34.929 42.24 36.888 ;
      RECT 42.234 34.883 42.286 36.842 ;
      RECT 42.28 34.837 42.332 36.796 ;
      RECT 42.326 34.791 42.378 36.75 ;
      RECT 42.372 34.745 42.424 36.704 ;
      RECT 42.418 34.699 42.47 36.658 ;
      RECT 42.464 34.653 42.516 36.612 ;
      RECT 42.51 34.607 42.562 36.566 ;
      RECT 42.556 34.561 42.608 36.52 ;
      RECT 42.602 34.515 42.654 36.474 ;
      RECT 42.648 34.469 42.7 36.428 ;
      RECT 42.694 34.423 42.746 36.382 ;
      RECT 42.74 34.377 42.792 36.336 ;
      RECT 42.786 34.331 42.838 36.29 ;
      RECT 42.832 34.285 42.884 36.244 ;
      RECT 42.878 34.239 42.93 36.198 ;
      RECT 42.924 34.193 42.976 36.152 ;
      RECT 42.97 34.147 43.022 36.106 ;
      RECT 43.016 34.101 43.068 36.06 ;
      RECT 43.062 34.055 43.114 36.014 ;
      RECT 43.108 34.009 43.16 35.968 ;
      RECT 43.154 33.963 43.206 35.922 ;
      RECT 43.2 33.917 43.252 35.876 ;
      RECT 43.246 33.871 43.298 35.83 ;
      RECT 43.292 33.825 43.344 35.784 ;
      RECT 43.338 33.779 43.39 35.738 ;
      RECT 43.384 33.733 43.436 35.692 ;
      RECT 43.43 33.687 43.482 35.646 ;
      RECT 43.476 33.641 43.528 35.6 ;
      RECT 43.522 33.595 43.574 35.554 ;
      RECT 43.568 33.549 43.62 35.508 ;
      RECT 43.614 33.503 43.666 35.462 ;
      RECT 43.66 33.457 43.712 35.416 ;
      RECT 43.706 33.411 43.758 35.37 ;
      RECT 43.752 33.365 43.804 35.324 ;
      RECT 43.798 33.319 43.85 35.278 ;
      RECT 43.844 33.273 43.896 35.232 ;
      RECT 43.89 33.227 43.942 35.186 ;
      RECT 43.936 33.181 43.988 35.14 ;
      RECT 43.982 33.135 44.034 35.094 ;
      RECT 44.028 33.089 44.08 35.048 ;
      RECT 44.074 33.043 44.126 35.002 ;
      RECT 44.12 32.997 44.172 34.956 ;
      RECT 44.166 32.951 44.218 34.91 ;
      RECT 44.212 32.905 44.264 34.864 ;
      RECT 44.258 32.859 44.31 34.818 ;
      RECT 44.304 32.813 44.356 34.772 ;
      RECT 44.35 32.767 44.402 34.726 ;
      RECT 44.396 32.721 44.448 34.68 ;
      RECT 44.442 32.675 44.494 34.634 ;
      RECT 44.488 32.629 44.54 34.588 ;
      RECT 44.534 32.583 44.586 34.542 ;
      RECT 44.58 32.537 44.632 34.496 ;
      RECT 44.626 32.491 44.678 34.45 ;
      RECT 44.672 32.445 44.724 34.404 ;
      RECT 44.718 32.399 44.77 34.358 ;
      RECT 44.764 32.353 44.816 34.312 ;
      RECT 44.81 32.307 44.862 34.266 ;
      RECT 44.856 32.261 44.908 34.22 ;
      RECT 44.902 32.215 44.954 34.174 ;
      RECT 44.948 32.169 45 34.128 ;
      RECT 44.994 32.123 45.046 34.082 ;
      RECT 45.04 32.077 45.092 34.036 ;
      RECT 45.086 32.031 45.138 33.99 ;
      RECT 45.132 31.985 45.184 33.944 ;
      RECT 45.178 31.939 45.23 33.898 ;
      RECT 45.224 31.893 45.276 33.852 ;
      RECT 45.27 31.847 45.322 33.806 ;
      RECT 45.316 31.801 45.368 33.76 ;
      RECT 45.362 31.755 45.414 33.714 ;
      RECT 45.408 31.709 45.46 33.668 ;
      RECT 45.454 31.663 45.506 33.622 ;
      RECT 45.5 31.617 45.552 33.576 ;
      RECT 45.546 31.571 45.598 33.53 ;
      RECT 45.592 31.525 45.644 33.484 ;
      RECT 45.638 31.479 45.69 33.438 ;
      RECT 45.684 31.433 45.736 33.392 ;
      RECT 45.73 31.387 45.782 33.346 ;
      RECT 45.776 31.341 45.828 33.3 ;
      RECT 45.822 31.295 45.874 33.254 ;
      RECT 45.868 31.249 45.92 33.208 ;
      RECT 45.914 31.203 45.966 33.162 ;
      RECT 45.96 31.157 46.012 33.116 ;
      RECT 46.006 31.111 46.058 33.07 ;
      RECT 46.052 31.065 46.104 33.024 ;
      RECT 46.098 31.019 46.15 32.978 ;
      RECT 46.144 30.973 46.196 32.932 ;
      RECT 46.19 30.927 46.242 32.886 ;
      RECT 46.236 30.881 46.288 32.84 ;
      RECT 46.282 30.835 46.334 32.794 ;
      RECT 46.328 30.789 46.38 32.748 ;
      RECT 46.374 30.743 46.426 32.702 ;
      RECT 46.42 30.697 46.472 32.656 ;
      RECT 46.466 30.651 46.518 32.61 ;
      RECT 46.512 30.605 46.564 32.564 ;
      RECT 46.558 30.559 46.61 32.518 ;
      RECT 46.604 30.513 46.656 32.472 ;
      RECT 46.65 30.467 46.702 32.426 ;
      RECT 46.696 30.421 46.748 32.38 ;
      RECT 46.742 30.375 46.794 32.334 ;
      RECT 46.788 30.329 46.84 32.288 ;
      RECT 46.834 30.283 46.886 32.242 ;
      RECT 46.88 30.237 46.932 32.196 ;
      RECT 46.926 30.191 46.978 32.15 ;
      RECT 46.972 30.145 47.024 32.104 ;
      RECT 47.018 30.099 47.07 32.058 ;
      RECT 47.064 30.053 47.116 32.012 ;
      RECT 47.11 30.007 47.162 31.966 ;
      RECT 47.156 29.961 47.208 31.92 ;
      RECT 47.202 29.915 47.254 31.874 ;
      RECT 47.248 29.869 47.3 31.828 ;
      RECT 47.294 29.823 47.346 31.782 ;
      RECT 47.34 29.777 47.392 31.736 ;
      RECT 47.386 29.731 47.438 31.69 ;
      RECT 47.432 29.685 47.484 31.644 ;
      RECT 47.478 29.639 47.53 31.598 ;
      RECT 47.524 29.593 47.576 31.552 ;
      RECT 47.57 29.547 47.622 31.506 ;
      RECT 47.616 29.501 47.668 31.46 ;
      RECT 47.662 29.455 47.714 31.414 ;
      RECT 47.708 29.409 47.76 31.368 ;
      RECT 47.754 29.363 47.806 31.322 ;
      RECT 47.8 29.317 47.852 31.276 ;
      RECT 47.846 29.271 47.898 31.23 ;
      RECT 47.892 29.225 47.944 31.184 ;
      RECT 47.938 29.179 47.99 31.138 ;
      RECT 47.984 29.133 48.036 31.092 ;
      RECT 48.03 29.087 48.082 31.046 ;
      RECT 48.076 29.041 48.128 31 ;
      RECT 48.122 28.995 48.174 30.954 ;
      RECT 48.168 28.949 48.22 30.908 ;
      RECT 48.214 28.903 48.266 30.862 ;
      RECT 48.26 28.857 48.312 30.816 ;
      RECT 48.306 28.811 48.358 30.77 ;
      RECT 48.352 28.765 48.404 30.724 ;
      RECT 48.398 28.719 48.45 30.678 ;
      RECT 48.444 28.673 48.496 30.632 ;
      RECT 48.49 28.627 48.542 30.586 ;
      RECT 48.536 28.581 48.588 30.54 ;
      RECT 48.582 28.535 48.634 30.494 ;
      RECT 48.628 28.489 48.68 30.448 ;
      RECT 48.674 28.443 48.726 30.402 ;
      RECT 48.72 28.397 48.772 30.356 ;
      RECT 48.766 28.351 48.818 30.31 ;
      RECT 48.812 28.305 48.864 30.264 ;
      RECT 48.858 28.259 48.91 30.218 ;
      RECT 48.904 28.213 48.956 30.172 ;
      RECT 48.95 28.167 49.002 30.126 ;
      RECT 48.996 28.121 49.048 30.08 ;
      RECT 49.042 28.075 49.094 30.034 ;
      RECT 49.088 28.029 49.14 29.988 ;
      RECT 49.134 27.983 49.186 29.942 ;
      RECT 49.18 27.937 49.232 29.896 ;
      RECT 49.226 27.891 49.278 29.85 ;
      RECT 49.272 27.845 49.324 29.804 ;
      RECT 49.318 27.799 49.37 29.758 ;
      RECT 49.364 27.753 49.416 29.712 ;
      RECT 49.41 27.707 49.462 29.666 ;
      RECT 49.456 27.661 49.508 29.62 ;
      RECT 49.502 27.615 49.554 29.574 ;
      RECT 49.548 27.569 49.6 29.528 ;
      RECT 49.594 27.523 49.646 29.482 ;
      RECT 49.64 27.477 49.692 29.436 ;
      RECT 49.686 27.431 49.738 29.39 ;
      RECT 49.732 27.385 49.784 29.344 ;
      RECT 49.778 27.339 49.83 29.298 ;
      RECT 49.824 27.293 49.876 29.252 ;
      RECT 49.87 27.247 49.922 29.206 ;
      RECT 49.916 27.201 49.968 29.16 ;
      RECT 49.962 27.155 50.014 29.114 ;
      RECT 50.008 27.109 50.06 29.068 ;
      RECT 50.054 27.063 50.106 29.022 ;
      RECT 50.1 27.017 50.152 28.976 ;
      RECT 50.146 26.971 50.198 28.93 ;
      RECT 50.192 26.925 50.244 28.884 ;
      RECT 50.238 26.879 50.29 28.838 ;
      RECT 50.284 26.833 50.336 28.792 ;
      RECT 50.33 26.787 50.382 28.746 ;
      RECT 50.376 26.741 50.428 28.7 ;
      RECT 50.422 26.695 50.474 28.654 ;
      RECT 50.468 26.649 50.52 28.608 ;
      RECT 50.514 26.603 50.566 28.562 ;
      RECT 50.56 26.557 50.612 28.516 ;
      RECT 50.606 26.511 50.658 28.47 ;
      RECT 50.652 26.465 50.704 28.424 ;
      RECT 50.698 26.419 50.75 28.378 ;
      RECT 50.744 26.373 50.796 28.332 ;
      RECT 50.79 26.327 50.842 28.286 ;
      RECT 50.836 26.281 50.888 28.24 ;
      RECT 50.882 26.235 50.934 28.194 ;
      RECT 50.928 26.189 50.98 28.148 ;
      RECT 50.974 26.143 51.026 28.102 ;
      RECT 51.02 26.097 51.072 28.056 ;
      RECT 51.066 26.051 51.118 28.01 ;
      RECT 51.112 26.005 51.164 27.964 ;
      RECT 51.158 25.959 51.21 27.918 ;
      RECT 51.204 25.913 51.256 27.872 ;
      RECT 51.25 25.867 51.302 27.826 ;
      RECT 51.296 25.821 51.348 27.78 ;
      RECT 51.342 25.775 51.394 27.734 ;
      RECT 51.388 25.729 51.44 27.688 ;
      RECT 51.434 25.683 51.486 27.642 ;
      RECT 51.48 25.637 51.532 27.596 ;
      RECT 51.526 25.591 51.578 27.55 ;
      RECT 51.572 25.545 51.624 27.504 ;
      RECT 51.618 25.499 51.67 27.458 ;
      RECT 51.664 25.453 51.716 27.412 ;
      RECT 51.71 25.407 51.762 27.366 ;
      RECT 51.756 25.361 51.808 27.32 ;
      RECT 51.802 25.315 51.854 27.274 ;
      RECT 51.848 25.269 51.9 27.228 ;
      RECT 51.894 25.223 51.946 27.182 ;
      RECT 51.94 25.177 51.992 27.136 ;
      RECT 51.986 25.131 52.038 27.09 ;
      RECT 52.032 25.085 52.084 27.044 ;
      RECT 52.078 25.039 52.13 26.998 ;
      RECT 52.124 24.993 52.176 26.952 ;
      RECT 52.17 24.947 52.222 26.906 ;
      RECT 52.216 24.901 52.268 26.86 ;
      RECT 52.262 24.855 52.314 26.814 ;
      RECT 52.308 24.809 52.36 26.768 ;
      RECT 52.354 24.763 52.406 26.722 ;
      RECT 52.4 24.717 52.452 26.676 ;
      RECT 52.446 24.671 52.498 26.63 ;
      RECT 52.492 24.625 52.544 26.584 ;
      RECT 52.538 24.579 52.59 26.538 ;
      RECT 52.584 24.533 52.636 26.492 ;
      RECT 52.63 24.487 52.682 26.446 ;
      RECT 52.676 24.441 52.728 26.4 ;
      RECT 52.722 24.395 52.774 26.354 ;
      RECT 52.768 24.349 52.82 26.308 ;
      RECT 52.814 24.303 52.866 26.262 ;
      RECT 52.86 24.257 52.912 26.216 ;
      RECT 52.906 24.211 52.958 26.17 ;
      RECT 52.952 24.165 53.004 26.124 ;
      RECT 52.998 24.119 53.05 26.078 ;
      RECT 53.044 24.073 53.096 26.032 ;
      RECT 53.09 24.027 53.142 25.986 ;
      RECT 53.136 23.981 53.188 25.94 ;
      RECT 53.182 23.935 53.234 25.894 ;
      RECT 53.228 23.889 53.28 25.848 ;
      RECT 53.274 23.843 53.326 25.802 ;
      RECT 53.32 23.797 53.372 25.756 ;
      RECT 53.366 23.751 53.418 25.71 ;
      RECT 53.412 23.705 53.464 25.664 ;
      RECT 53.458 23.659 53.51 25.618 ;
      RECT 53.504 23.613 53.556 25.572 ;
      RECT 53.55 23.567 53.602 25.526 ;
      RECT 53.596 23.521 53.648 25.48 ;
      RECT 53.642 23.475 53.694 25.434 ;
      RECT 53.688 23.429 53.74 25.388 ;
      RECT 53.734 23.383 53.786 25.342 ;
      RECT 53.78 23.337 53.832 25.296 ;
      RECT 53.826 23.291 53.878 25.25 ;
      RECT 53.872 23.245 53.924 25.204 ;
      RECT 53.918 23.199 53.97 25.158 ;
      RECT 53.964 23.153 54.016 25.112 ;
      RECT 54.01 23.107 54.062 25.066 ;
      RECT 54.056 23.061 54.108 25.02 ;
      RECT 54.102 23.015 54.154 24.974 ;
      RECT 54.148 22.969 54.2 24.928 ;
      RECT 54.194 22.923 54.246 24.882 ;
      RECT 54.24 22.877 54.292 24.836 ;
      RECT 54.286 22.831 54.338 24.79 ;
      RECT 54.332 22.785 54.384 24.744 ;
      RECT 54.378 22.739 54.43 24.698 ;
      RECT 54.424 22.693 54.476 24.652 ;
      RECT 54.47 22.647 54.522 24.606 ;
      RECT 54.516 22.601 54.568 24.56 ;
      RECT 54.562 22.555 54.614 24.514 ;
      RECT 54.608 22.509 54.66 24.468 ;
      RECT 54.654 22.463 54.706 24.422 ;
      RECT 54.7 22.417 54.752 24.376 ;
      RECT 54.746 22.371 54.798 24.33 ;
      RECT 54.792 22.325 54.844 24.284 ;
      RECT 54.838 22.279 54.89 24.238 ;
      RECT 54.884 22.233 54.936 24.192 ;
      RECT 54.93 22.187 54.982 24.146 ;
      RECT 54.976 22.141 55.028 24.1 ;
      RECT 55.022 22.095 55.074 24.054 ;
      RECT 55.068 22.049 55.12 24.008 ;
      RECT 55.114 22.003 55.166 23.962 ;
      RECT 55.16 21.957 55.212 23.916 ;
      RECT 55.206 21.911 55.258 23.87 ;
      RECT 55.252 21.865 55.304 23.824 ;
      RECT 55.298 21.819 55.35 23.778 ;
      RECT 55.344 21.773 55.396 23.732 ;
      RECT 55.39 21.727 55.442 23.686 ;
      RECT 55.436 21.681 55.488 23.64 ;
      RECT 55.482 21.635 55.534 23.594 ;
      RECT 55.528 21.589 55.58 23.548 ;
      RECT 55.574 21.543 55.626 23.502 ;
      RECT 55.62 21.497 55.672 23.456 ;
      RECT 55.666 21.451 55.718 23.41 ;
      RECT 55.712 21.405 55.764 23.364 ;
      RECT 55.758 21.359 55.81 23.318 ;
      RECT 55.804 21.313 55.856 23.272 ;
      RECT 55.85 21.267 55.902 23.226 ;
      RECT 55.896 21.221 55.948 23.18 ;
      RECT 55.942 21.175 55.994 23.134 ;
      RECT 55.988 21.129 56.04 23.088 ;
      RECT 56.034 21.083 56.086 23.042 ;
      RECT 56.08 21.037 56.132 22.996 ;
      RECT 56.126 20.991 56.178 22.95 ;
      RECT 56.172 20.945 56.224 22.904 ;
      RECT 56.218 20.899 56.27 22.858 ;
      RECT 56.264 20.853 56.316 22.812 ;
      RECT 56.31 20.813 56.362 22.766 ;
      RECT 56.345 20.772 56.408 22.72 ;
      RECT 56.391 20.726 56.454 22.674 ;
      RECT 56.437 20.68 56.5 22.628 ;
      RECT 56.483 20.634 56.546 22.582 ;
      RECT 56.529 20.588 56.592 22.536 ;
      RECT 56.575 20.542 56.638 22.49 ;
      RECT 56.621 20.496 56.684 22.444 ;
      RECT 56.667 20.45 56.73 22.398 ;
      RECT 56.713 20.404 56.776 22.352 ;
      RECT 56.759 20.358 56.822 22.306 ;
      RECT 56.805 20.312 56.868 22.26 ;
      RECT 56.851 20.266 56.914 22.214 ;
      RECT 56.897 20.22 56.96 22.168 ;
      RECT 56.943 20.174 57.006 22.122 ;
      RECT 56.989 20.128 57.052 22.076 ;
      RECT 57.035 20.082 57.098 22.03 ;
      RECT 57.081 20.036 57.144 21.984 ;
      RECT 57.127 19.99 57.19 21.938 ;
      RECT 57.173 19.944 57.236 21.892 ;
      RECT 57.219 19.898 57.282 21.846 ;
      RECT 57.265 19.852 57.328 21.8 ;
      RECT 57.311 19.806 57.374 21.754 ;
      RECT 57.357 19.76 57.42 21.708 ;
      RECT 57.403 19.714 57.466 21.662 ;
      RECT 57.449 19.668 57.512 21.616 ;
      RECT 57.495 19.622 57.558 21.57 ;
      RECT 57.541 19.576 57.604 21.524 ;
      RECT 57.587 19.53 57.65 21.478 ;
      RECT 57.633 19.484 57.696 21.432 ;
      RECT 57.679 19.438 57.742 21.386 ;
      RECT 57.725 19.392 57.788 21.34 ;
      RECT 57.771 19.346 57.834 21.294 ;
      RECT 57.817 19.3 57.88 21.248 ;
      RECT 57.863 19.254 57.926 21.202 ;
      RECT 57.909 19.208 57.972 21.156 ;
      RECT 57.955 19.162 58.018 21.11 ;
      RECT 58.001 19.116 58.064 21.064 ;
      RECT 58.047 19.07 58.11 21.018 ;
      RECT 58.093 19.024 58.156 20.972 ;
      RECT 58.139 18.978 58.202 20.926 ;
      RECT 58.185 18.932 58.248 20.88 ;
      RECT 58.231 18.886 58.294 20.834 ;
      RECT 58.277 18.84 58.34 20.788 ;
      RECT 58.323 18.794 58.386 20.742 ;
      RECT 58.369 18.748 58.432 20.696 ;
      RECT 58.415 18.702 58.478 20.65 ;
      RECT 58.461 18.656 58.524 20.604 ;
      RECT 58.507 18.61 58.57 20.558 ;
      RECT 58.553 18.564 58.616 20.512 ;
      RECT 58.599 18.518 58.662 20.466 ;
      RECT 58.645 18.472 58.708 20.42 ;
      RECT 58.691 18.426 58.754 20.374 ;
      RECT 58.737 18.38 58.8 20.328 ;
      RECT 58.783 18.334 58.846 20.282 ;
      RECT 58.829 18.288 58.892 20.236 ;
      RECT 58.875 18.242 58.938 20.19 ;
      RECT 58.921 18.196 58.984 20.144 ;
      RECT 58.967 18.15 59.03 20.098 ;
      RECT 59.013 18.104 59.076 20.052 ;
      RECT 59.059 18.058 59.122 20.006 ;
      RECT 59.105 18.012 59.168 19.96 ;
      RECT 59.151 17.966 59.214 19.914 ;
      RECT 59.197 17.92 59.26 19.868 ;
      RECT 59.243 17.874 59.306 19.822 ;
      RECT 59.289 17.828 59.352 19.776 ;
      RECT 59.335 17.782 59.398 19.73 ;
      RECT 59.381 17.736 59.444 19.684 ;
      RECT 59.427 17.69 59.49 19.638 ;
      RECT 59.473 17.644 59.536 19.592 ;
      RECT 59.519 17.598 59.582 19.546 ;
      RECT 59.565 17.552 59.628 19.5 ;
      RECT 59.611 17.506 59.674 19.454 ;
      RECT 59.657 17.46 59.72 19.408 ;
      RECT 59.703 17.414 59.766 19.362 ;
      RECT 59.749 17.368 59.812 19.316 ;
      RECT 59.795 17.322 59.858 19.27 ;
      RECT 59.841 17.276 59.904 19.224 ;
      RECT 59.887 17.23 59.95 19.178 ;
      RECT 59.933 17.184 59.996 19.132 ;
      RECT 59.979 17.138 60.042 19.086 ;
      RECT 60.025 17.092 60.088 19.04 ;
      RECT 60.071 17.046 60.134 18.994 ;
      RECT 60.117 17 60.18 18.948 ;
      RECT 60.163 16.954 60.226 18.902 ;
      RECT 60.209 16.908 60.272 18.856 ;
      RECT 60.255 16.862 60.318 18.81 ;
      RECT 60.301 16.816 60.364 18.764 ;
      RECT 60.347 16.77 60.41 18.718 ;
      RECT 60.393 16.724 60.456 18.672 ;
      RECT 60.439 16.678 60.502 18.626 ;
      RECT 60.485 16.632 60.548 18.58 ;
      RECT 60.531 16.586 60.594 18.534 ;
      RECT 60.577 16.54 60.64 18.488 ;
      RECT 60.623 16.494 60.686 18.442 ;
      RECT 60.669 16.448 60.732 18.396 ;
      RECT 60.715 16.402 60.778 18.35 ;
      RECT 60.761 16.356 60.824 18.304 ;
      RECT 60.807 16.31 60.87 18.258 ;
      RECT 60.853 16.264 60.916 18.212 ;
      RECT 60.899 16.218 60.962 18.166 ;
      RECT 60.945 16.172 61.008 18.12 ;
      RECT 60.991 16.126 61.054 18.074 ;
      RECT 61.037 16.08 61.1 18.028 ;
      RECT 61.083 16.034 61.146 17.982 ;
      RECT 61.129 15.988 61.192 17.936 ;
      RECT 61.175 15.942 61.238 17.89 ;
      RECT 61.221 15.896 61.284 17.844 ;
      RECT 61.267 15.852 61.33 17.798 ;
      RECT 61.31 15.83 61.376 17.752 ;
      RECT 61.31 15.83 61.422 17.706 ;
      RECT 61.31 15.83 61.468 17.66 ;
      RECT 61.31 15.83 61.514 17.614 ;
      RECT 61.31 15.83 61.56 17.568 ;
      RECT 61.31 15.83 61.606 17.522 ;
      RECT 61.31 15.83 61.652 17.476 ;
      RECT 61.31 15.83 61.698 17.43 ;
      RECT 61.31 15.83 61.744 17.384 ;
      RECT 61.31 15.83 61.79 17.338 ;
      RECT 61.31 15.83 61.836 17.292 ;
      RECT 61.31 15.83 61.882 17.246 ;
      RECT 61.31 15.83 61.928 17.2 ;
      RECT 61.31 15.83 61.974 17.154 ;
      RECT 61.31 15.83 62.02 17.108 ;
      RECT 61.31 15.83 62.066 17.062 ;
      RECT 61.31 15.83 62.112 17.016 ;
      RECT 61.31 15.83 62.158 16.97 ;
      RECT 61.31 15.83 62.204 16.924 ;
      RECT 61.31 15.83 62.25 16.878 ;
      RECT 61.31 15.83 62.296 16.832 ;
      RECT 61.31 15.83 62.342 16.786 ;
      RECT 61.31 15.83 62.388 16.74 ;
      RECT 61.31 15.83 62.434 16.694 ;
      RECT 61.31 15.83 110 16.67 ;
      RECT 29.33 68.037 30.17 110 ;
      RECT 29.33 68.037 30.216 69.162 ;
      RECT 29.33 68.037 30.262 69.116 ;
      RECT 29.33 68.037 30.308 69.07 ;
      RECT 29.33 68.037 30.354 69.024 ;
      RECT 29.33 68.037 30.4 68.978 ;
      RECT 29.33 68.037 30.446 68.932 ;
      RECT 29.33 68.037 30.492 68.886 ;
      RECT 29.33 68.037 30.538 68.84 ;
      RECT 29.33 68.037 30.584 68.794 ;
      RECT 29.33 68.037 30.63 68.748 ;
      RECT 29.33 68.037 30.676 68.702 ;
      RECT 29.33 68.037 30.722 68.656 ;
      RECT 29.33 68.037 30.768 68.61 ;
      RECT 29.33 68.037 30.814 68.564 ;
      RECT 29.33 68.037 30.86 68.518 ;
      RECT 29.33 68.037 30.906 68.472 ;
      RECT 29.33 68.037 30.952 68.426 ;
      RECT 29.33 68.037 30.998 68.38 ;
      RECT 29.33 68.037 31.044 68.334 ;
      RECT 29.33 68.037 31.09 68.288 ;
      RECT 29.33 68.037 31.136 68.242 ;
      RECT 29.33 68.037 31.182 68.196 ;
      RECT 29.33 68.037 31.228 68.15 ;
      RECT 29.33 68.037 31.274 68.104 ;
      RECT 29.376 67.991 31.32 68.058 ;
      RECT 29.422 67.945 31.366 68.012 ;
      RECT 29.468 67.899 31.412 67.966 ;
      RECT 29.514 67.853 31.458 67.92 ;
      RECT 29.56 67.807 31.504 67.874 ;
      RECT 29.606 67.761 31.55 67.828 ;
      RECT 29.652 67.715 31.596 67.782 ;
      RECT 29.698 67.669 31.642 67.736 ;
      RECT 29.744 67.623 31.688 67.69 ;
      RECT 29.79 67.577 31.734 67.644 ;
      RECT 29.836 67.531 31.78 67.598 ;
      RECT 29.882 67.485 31.826 67.552 ;
      RECT 29.928 67.439 31.872 67.506 ;
      RECT 29.974 67.393 31.918 67.46 ;
      RECT 30.02 67.347 31.964 67.414 ;
      RECT 30.066 67.301 32.01 67.368 ;
      RECT 30.112 67.255 32.056 67.322 ;
      RECT 30.158 67.209 32.102 67.276 ;
      RECT 30.204 67.163 32.148 67.23 ;
      RECT 30.25 67.117 32.194 67.184 ;
      RECT 30.296 67.071 32.24 67.138 ;
      RECT 30.342 67.025 32.286 67.092 ;
      RECT 30.388 66.979 32.332 67.046 ;
      RECT 30.434 66.933 32.378 67 ;
      RECT 30.48 66.887 32.424 66.954 ;
      RECT 30.526 66.841 32.47 66.908 ;
      RECT 30.572 66.795 32.516 66.862 ;
      RECT 30.618 66.749 32.562 66.816 ;
      RECT 30.664 66.703 32.608 66.77 ;
      RECT 30.71 66.657 32.654 66.724 ;
      RECT 30.756 66.611 32.7 66.678 ;
      RECT 30.802 66.565 32.746 66.632 ;
      RECT 30.848 66.519 32.792 66.586 ;
      RECT 30.894 66.473 32.838 66.54 ;
      RECT 30.94 66.427 32.884 66.494 ;
      RECT 30.986 66.381 32.93 66.448 ;
      RECT 31.032 66.335 32.976 66.402 ;
      RECT 31.078 66.289 33.022 66.356 ;
      RECT 31.124 66.243 33.068 66.31 ;
      RECT 31.17 66.197 33.114 66.264 ;
      RECT 31.216 66.151 33.16 66.218 ;
      RECT 31.262 66.105 33.206 66.172 ;
      RECT 31.308 66.059 33.252 66.126 ;
      RECT 31.354 66.013 33.298 66.08 ;
      RECT 31.4 65.967 33.344 66.034 ;
      RECT 31.446 65.921 33.39 65.988 ;
      RECT 31.492 65.875 33.436 65.942 ;
      RECT 31.538 65.829 33.482 65.896 ;
      RECT 31.584 65.783 33.528 65.85 ;
      RECT 31.63 65.737 33.574 65.804 ;
      RECT 31.676 65.691 33.62 65.758 ;
      RECT 31.722 65.645 33.666 65.712 ;
      RECT 31.768 65.599 33.712 65.666 ;
      RECT 31.814 65.553 33.758 65.62 ;
      RECT 31.86 65.507 33.804 65.574 ;
      RECT 31.906 65.461 33.85 65.528 ;
      RECT 31.952 65.415 33.896 65.482 ;
      RECT 31.998 65.369 33.942 65.436 ;
      RECT 32.044 65.323 33.988 65.39 ;
      RECT 32.09 65.277 34.034 65.344 ;
      RECT 32.136 65.231 34.08 65.298 ;
      RECT 32.182 65.185 34.126 65.252 ;
      RECT 32.228 65.139 34.172 65.206 ;
      RECT 32.274 65.093 34.218 65.16 ;
      RECT 32.32 65.047 34.264 65.114 ;
      RECT 32.366 65.001 34.31 65.068 ;
      RECT 32.412 64.955 34.356 65.022 ;
      RECT 32.458 64.909 34.402 64.976 ;
      RECT 32.504 64.863 34.448 64.93 ;
      RECT 32.55 64.817 34.494 64.884 ;
      RECT 32.596 64.771 34.54 64.838 ;
      RECT 32.642 64.725 34.586 64.792 ;
      RECT 32.688 64.679 34.632 64.746 ;
      RECT 32.734 64.633 34.678 64.7 ;
      RECT 32.78 64.587 34.724 64.654 ;
      RECT 32.826 64.541 34.77 64.608 ;
      RECT 32.872 64.495 34.816 64.562 ;
      RECT 32.918 64.449 34.862 64.516 ;
      RECT 32.964 64.403 34.908 64.47 ;
      RECT 33.01 64.357 34.954 64.424 ;
      RECT 33.056 64.311 35 64.378 ;
      RECT 33.102 64.265 35.046 64.332 ;
      RECT 33.148 64.219 35.092 64.286 ;
      RECT 33.194 64.173 35.138 64.24 ;
      RECT 33.24 64.127 35.184 64.194 ;
      RECT 33.286 64.081 35.23 64.148 ;
      RECT 33.332 64.035 35.276 64.102 ;
      RECT 33.378 63.989 35.322 64.056 ;
      RECT 33.424 63.943 35.368 64.01 ;
      RECT 33.47 63.897 35.414 63.964 ;
      RECT 33.516 63.851 35.46 63.918 ;
      RECT 33.562 63.805 35.506 63.872 ;
      RECT 33.608 63.759 35.552 63.826 ;
      RECT 33.654 63.713 35.598 63.78 ;
      RECT 33.7 63.667 35.644 63.734 ;
      RECT 33.746 63.621 35.69 63.688 ;
      RECT 33.792 63.575 35.736 63.642 ;
      RECT 33.838 63.529 35.782 63.596 ;
      RECT 33.884 63.483 35.828 63.55 ;
      RECT 33.93 63.437 35.874 63.504 ;
      RECT 33.976 63.391 35.92 63.458 ;
      RECT 34.022 63.345 35.966 63.412 ;
      RECT 34.068 63.299 36.012 63.366 ;
      RECT 34.114 63.253 36.058 63.32 ;
      RECT 34.16 63.207 36.104 63.274 ;
      RECT 34.206 63.161 36.15 63.228 ;
      RECT 34.252 63.115 36.196 63.182 ;
      RECT 34.298 63.069 36.242 63.136 ;
      RECT 34.344 63.023 36.288 63.09 ;
      RECT 34.39 62.977 36.334 63.044 ;
      RECT 34.436 62.931 36.38 62.998 ;
      RECT 34.482 62.885 36.426 62.952 ;
      RECT 34.528 62.839 36.472 62.906 ;
      RECT 34.574 62.793 36.518 62.86 ;
      RECT 34.62 62.747 36.564 62.814 ;
      RECT 34.666 62.701 36.61 62.768 ;
      RECT 34.712 62.655 36.656 62.722 ;
      RECT 34.758 62.609 36.702 62.676 ;
      RECT 34.804 62.563 36.748 62.63 ;
      RECT 34.85 62.517 36.794 62.584 ;
      RECT 34.896 62.471 36.84 62.538 ;
      RECT 34.942 62.425 36.886 62.492 ;
      RECT 34.988 62.379 36.932 62.446 ;
      RECT 35.034 62.333 36.978 62.4 ;
      RECT 35.08 62.287 37.024 62.354 ;
      RECT 35.126 62.241 37.07 62.308 ;
      RECT 35.172 62.195 37.116 62.262 ;
      RECT 35.218 62.149 37.162 62.216 ;
      RECT 35.264 62.103 37.208 62.17 ;
      RECT 35.31 62.057 37.254 62.124 ;
      RECT 35.356 62.011 37.3 62.078 ;
      RECT 35.402 61.965 37.346 62.032 ;
      RECT 35.448 61.919 37.392 61.986 ;
      RECT 35.494 61.873 37.438 61.94 ;
      RECT 35.54 61.827 37.484 61.894 ;
      RECT 35.586 61.781 37.53 61.848 ;
      RECT 35.632 61.735 37.576 61.802 ;
      RECT 35.678 61.689 37.622 61.756 ;
      RECT 35.724 61.643 37.668 61.71 ;
      RECT 35.77 61.597 37.714 61.664 ;
      RECT 35.816 61.551 37.76 61.618 ;
      RECT 35.862 61.505 37.806 61.572 ;
      RECT 35.908 61.459 37.852 61.526 ;
      RECT 35.954 61.413 37.898 61.48 ;
      RECT 36 61.367 37.944 61.434 ;
      RECT 36.046 61.321 37.99 61.388 ;
      RECT 36.092 61.275 38.036 61.342 ;
      RECT 36.138 61.229 38.082 61.296 ;
      RECT 36.184 61.183 38.128 61.25 ;
      RECT 36.23 61.137 38.174 61.204 ;
      RECT 36.276 61.091 38.22 61.158 ;
      RECT 36.322 61.045 38.266 61.112 ;
      RECT 36.368 60.999 38.312 61.066 ;
      RECT 36.414 60.953 38.358 61.02 ;
      RECT 36.46 60.907 38.404 60.974 ;
      RECT 36.506 60.861 38.45 60.928 ;
      RECT 36.552 60.815 38.496 60.882 ;
      RECT 36.598 60.769 38.542 60.836 ;
      RECT 36.644 60.723 38.588 60.79 ;
      RECT 36.69 60.677 38.634 60.744 ;
      RECT 36.736 60.631 38.68 60.698 ;
      RECT 36.782 60.585 38.726 60.652 ;
      RECT 36.828 60.539 38.772 60.606 ;
      RECT 36.874 60.493 38.818 60.56 ;
      RECT 36.92 60.447 38.864 60.514 ;
      RECT 36.966 60.401 38.91 60.468 ;
      RECT 37.012 60.355 38.956 60.422 ;
      RECT 37.058 60.309 39.002 60.376 ;
      RECT 37.104 60.263 39.048 60.33 ;
      RECT 37.15 60.217 39.094 60.284 ;
      RECT 37.196 60.171 39.14 60.238 ;
      RECT 37.242 60.125 39.186 60.192 ;
      RECT 37.288 60.079 39.232 60.146 ;
      RECT 37.334 60.033 39.278 60.1 ;
      RECT 37.38 59.987 39.324 60.054 ;
      RECT 37.426 59.941 39.37 60.008 ;
      RECT 37.472 59.895 39.416 59.962 ;
      RECT 37.518 59.849 39.462 59.916 ;
      RECT 37.564 59.803 39.508 59.87 ;
      RECT 37.61 59.757 39.554 59.824 ;
      RECT 37.656 59.711 39.6 59.778 ;
      RECT 37.702 59.665 39.646 59.732 ;
      RECT 37.748 59.619 39.692 59.686 ;
      RECT 37.794 59.573 39.738 59.64 ;
      RECT 37.84 59.527 39.784 59.594 ;
      RECT 37.886 59.481 39.83 59.548 ;
      RECT 37.932 59.435 39.876 59.502 ;
      RECT 37.978 59.389 39.922 59.456 ;
      RECT 38.024 59.343 39.968 59.41 ;
      RECT 38.07 59.297 40.014 59.364 ;
      RECT 38.116 59.251 40.06 59.318 ;
      RECT 38.162 59.205 40.106 59.272 ;
      RECT 38.208 59.159 40.152 59.226 ;
      RECT 38.254 59.113 40.198 59.18 ;
      RECT 38.3 59.067 40.244 59.134 ;
      RECT 38.346 59.021 40.29 59.088 ;
      RECT 38.392 58.975 40.336 59.042 ;
      RECT 38.438 58.929 40.382 58.996 ;
      RECT 38.484 58.883 40.428 58.95 ;
      RECT 38.53 58.837 40.474 58.904 ;
      RECT 38.576 58.791 40.52 58.858 ;
      RECT 38.622 58.745 40.566 58.812 ;
      RECT 38.668 58.699 40.612 58.766 ;
      RECT 38.714 58.653 40.658 58.72 ;
      RECT 38.76 58.607 40.704 58.674 ;
      RECT 38.806 58.561 40.75 58.628 ;
      RECT 38.852 58.515 40.796 58.582 ;
      RECT 38.898 58.469 40.842 58.536 ;
      RECT 38.944 58.423 40.888 58.49 ;
      RECT 38.99 58.377 40.934 58.444 ;
      RECT 39.036 58.331 40.98 58.398 ;
      RECT 39.082 58.285 41.026 58.352 ;
      RECT 39.128 58.239 41.072 58.306 ;
      RECT 39.174 58.193 41.118 58.26 ;
      RECT 39.22 58.147 41.164 58.214 ;
      RECT 39.266 58.101 41.21 58.168 ;
      RECT 39.312 58.055 41.256 58.122 ;
      RECT 39.358 58.009 41.302 58.076 ;
      RECT 39.404 57.963 41.348 58.03 ;
      RECT 39.45 57.917 41.394 57.984 ;
      RECT 39.496 57.871 41.44 57.938 ;
      RECT 39.542 57.825 41.486 57.892 ;
      RECT 39.588 57.779 41.532 57.846 ;
      RECT 39.634 57.733 41.578 57.8 ;
      RECT 39.68 57.687 41.624 57.754 ;
      RECT 39.726 57.641 41.67 57.708 ;
      RECT 39.772 57.595 41.716 57.662 ;
      RECT 39.818 57.549 41.762 57.616 ;
      RECT 39.864 57.503 41.808 57.57 ;
      RECT 39.91 57.457 41.854 57.524 ;
      RECT 39.956 57.411 41.9 57.478 ;
      RECT 40.002 57.365 41.946 57.432 ;
      RECT 40.048 57.319 41.992 57.386 ;
      RECT 40.094 57.273 42.038 57.34 ;
      RECT 40.14 57.227 42.084 57.294 ;
      RECT 40.186 57.181 42.13 57.248 ;
      RECT 40.232 57.135 42.17 57.205 ;
      RECT 40.278 57.089 42.216 57.162 ;
      RECT 40.324 57.043 42.262 57.116 ;
      RECT 40.37 56.997 42.308 57.07 ;
      RECT 40.416 56.951 42.354 57.024 ;
      RECT 40.462 56.905 42.4 56.978 ;
      RECT 40.508 56.859 42.446 56.932 ;
      RECT 40.554 56.813 42.492 56.886 ;
      RECT 40.6 56.767 42.538 56.84 ;
      RECT 40.646 56.721 42.584 56.794 ;
      RECT 40.692 56.675 42.63 56.748 ;
      RECT 40.738 56.629 42.676 56.702 ;
      RECT 40.784 56.583 42.722 56.656 ;
      RECT 40.83 56.537 42.768 56.61 ;
      RECT 40.876 56.491 42.814 56.564 ;
      RECT 40.922 56.445 42.86 56.518 ;
      RECT 40.968 56.399 42.906 56.472 ;
      RECT 41.014 56.353 42.952 56.426 ;
      RECT 41.06 56.307 42.998 56.38 ;
      RECT 41.106 56.261 43.044 56.334 ;
      RECT 41.152 56.215 43.09 56.288 ;
      RECT 41.198 56.169 43.136 56.242 ;
      RECT 41.244 56.123 43.182 56.196 ;
      RECT 41.29 56.077 43.228 56.15 ;
      RECT 41.336 56.031 43.274 56.104 ;
      RECT 41.382 55.985 43.32 56.058 ;
      RECT 41.428 55.939 43.366 56.012 ;
      RECT 41.474 55.893 43.412 55.966 ;
      RECT 41.52 55.847 43.458 55.92 ;
      RECT 41.566 55.801 43.504 55.874 ;
      RECT 41.612 55.755 43.55 55.828 ;
      RECT 41.658 55.709 43.596 55.782 ;
      RECT 41.704 55.663 43.642 55.736 ;
      RECT 41.75 55.617 43.688 55.69 ;
      RECT 41.796 55.571 43.734 55.644 ;
      RECT 41.842 55.525 43.78 55.598 ;
      RECT 41.888 55.479 43.826 55.552 ;
      RECT 41.934 55.433 43.872 55.506 ;
      RECT 41.98 55.387 43.918 55.46 ;
      RECT 42.026 55.341 43.964 55.414 ;
      RECT 42.072 55.295 44.01 55.368 ;
      RECT 42.118 55.249 44.056 55.322 ;
      RECT 42.164 55.203 44.102 55.276 ;
      RECT 42.21 55.157 44.148 55.23 ;
      RECT 42.256 55.111 44.194 55.184 ;
      RECT 42.302 55.065 44.24 55.138 ;
      RECT 42.348 55.019 44.286 55.092 ;
      RECT 42.394 54.973 44.332 55.046 ;
      RECT 42.44 54.927 44.378 55 ;
      RECT 42.486 54.881 44.424 54.954 ;
      RECT 42.532 54.835 44.47 54.908 ;
      RECT 42.578 54.789 44.516 54.862 ;
      RECT 42.624 54.743 44.562 54.816 ;
      RECT 42.67 54.697 44.608 54.77 ;
      RECT 42.716 54.651 44.654 54.724 ;
      RECT 42.762 54.605 44.7 54.678 ;
      RECT 42.808 54.559 44.746 54.632 ;
      RECT 42.854 54.513 44.792 54.586 ;
      RECT 42.9 54.467 44.838 54.54 ;
      RECT 42.946 54.421 44.884 54.494 ;
      RECT 42.992 54.375 44.93 54.448 ;
      RECT 43.038 54.329 44.976 54.402 ;
      RECT 43.084 54.283 45.022 54.356 ;
      RECT 43.13 54.237 45.068 54.31 ;
      RECT 43.176 54.191 45.114 54.264 ;
      RECT 43.222 54.145 45.16 54.218 ;
      RECT 43.268 54.099 45.206 54.172 ;
      RECT 43.314 54.053 45.252 54.126 ;
      RECT 43.36 54.007 45.298 54.08 ;
      RECT 43.406 53.961 45.344 54.034 ;
      RECT 43.452 53.915 45.39 53.988 ;
      RECT 43.498 53.869 45.436 53.942 ;
      RECT 43.544 53.823 45.482 53.896 ;
      RECT 43.59 53.777 45.528 53.85 ;
      RECT 43.636 53.731 45.574 53.804 ;
      RECT 43.682 53.685 45.62 53.758 ;
      RECT 43.728 53.639 45.666 53.712 ;
      RECT 43.774 53.593 45.712 53.666 ;
      RECT 43.82 53.547 45.758 53.62 ;
      RECT 43.866 53.501 45.804 53.574 ;
      RECT 43.912 53.455 45.85 53.528 ;
      RECT 43.958 53.409 45.896 53.482 ;
      RECT 44.004 53.363 45.942 53.436 ;
      RECT 44.05 53.317 45.988 53.39 ;
      RECT 44.096 53.271 46.034 53.344 ;
      RECT 44.142 53.225 46.08 53.298 ;
      RECT 44.188 53.179 46.126 53.252 ;
      RECT 44.234 53.133 46.172 53.206 ;
      RECT 44.28 53.087 46.218 53.16 ;
      RECT 44.326 53.041 46.264 53.114 ;
      RECT 44.372 52.995 46.31 53.068 ;
      RECT 44.418 52.949 46.356 53.022 ;
      RECT 44.464 52.903 46.402 52.976 ;
      RECT 44.51 52.857 46.448 52.93 ;
      RECT 44.556 52.811 46.494 52.884 ;
      RECT 44.602 52.765 46.54 52.838 ;
      RECT 44.648 52.719 46.586 52.792 ;
      RECT 44.694 52.673 46.632 52.746 ;
      RECT 44.74 52.627 46.678 52.7 ;
      RECT 44.786 52.581 46.724 52.654 ;
      RECT 44.832 52.535 46.77 52.608 ;
      RECT 44.878 52.489 46.816 52.562 ;
      RECT 44.924 52.443 46.862 52.516 ;
      RECT 44.97 52.397 46.908 52.47 ;
      RECT 45.016 52.351 46.954 52.424 ;
      RECT 45.062 52.305 47 52.378 ;
      RECT 45.108 52.259 47.046 52.332 ;
      RECT 45.154 52.213 47.092 52.286 ;
      RECT 45.2 52.167 47.138 52.24 ;
      RECT 45.246 52.121 47.184 52.194 ;
      RECT 45.292 52.075 47.23 52.148 ;
      RECT 45.338 52.029 47.276 52.102 ;
      RECT 45.384 51.983 47.322 52.056 ;
      RECT 45.43 51.937 47.368 52.01 ;
      RECT 45.476 51.891 47.414 51.964 ;
      RECT 45.522 51.845 47.46 51.918 ;
      RECT 45.568 51.799 47.506 51.872 ;
      RECT 45.614 51.753 47.552 51.826 ;
      RECT 45.66 51.707 47.598 51.78 ;
      RECT 45.706 51.661 47.644 51.734 ;
      RECT 45.752 51.615 47.69 51.688 ;
      RECT 45.798 51.569 47.736 51.642 ;
      RECT 45.844 51.523 47.782 51.596 ;
      RECT 45.89 51.477 47.828 51.55 ;
      RECT 45.936 51.431 47.874 51.504 ;
      RECT 45.982 51.385 47.92 51.458 ;
      RECT 46.028 51.339 47.966 51.412 ;
      RECT 46.074 51.293 48.012 51.366 ;
      RECT 46.12 51.247 48.058 51.32 ;
      RECT 46.166 51.201 48.104 51.274 ;
      RECT 46.212 51.155 48.15 51.228 ;
      RECT 46.258 51.109 48.196 51.182 ;
      RECT 46.304 51.063 48.242 51.136 ;
      RECT 46.35 51.017 48.288 51.09 ;
      RECT 46.396 50.971 48.334 51.044 ;
      RECT 46.442 50.925 48.38 50.998 ;
      RECT 46.488 50.879 48.426 50.952 ;
      RECT 46.534 50.833 48.472 50.906 ;
      RECT 46.58 50.787 48.518 50.86 ;
      RECT 46.626 50.741 48.564 50.814 ;
      RECT 46.672 50.695 48.61 50.768 ;
      RECT 46.718 50.649 48.656 50.722 ;
      RECT 46.764 50.603 48.702 50.676 ;
      RECT 46.81 50.557 48.748 50.63 ;
      RECT 46.856 50.511 48.794 50.584 ;
      RECT 46.902 50.465 48.84 50.538 ;
      RECT 46.948 50.419 48.886 50.492 ;
      RECT 46.994 50.373 48.932 50.446 ;
      RECT 47.04 50.327 48.978 50.4 ;
      RECT 47.086 50.281 49.024 50.354 ;
      RECT 47.132 50.235 49.07 50.308 ;
      RECT 47.178 50.189 49.116 50.262 ;
      RECT 47.224 50.143 49.162 50.216 ;
      RECT 47.27 50.097 49.208 50.17 ;
      RECT 47.316 50.051 49.254 50.124 ;
      RECT 47.362 50.005 49.3 50.078 ;
      RECT 47.408 49.959 49.346 50.032 ;
      RECT 47.454 49.913 49.392 49.986 ;
      RECT 47.5 49.867 49.438 49.94 ;
      RECT 47.546 49.821 49.484 49.894 ;
      RECT 47.592 49.775 49.53 49.848 ;
      RECT 47.638 49.729 49.576 49.802 ;
      RECT 47.684 49.683 49.622 49.756 ;
      RECT 47.73 49.637 49.668 49.71 ;
      RECT 47.776 49.591 49.714 49.664 ;
      RECT 47.822 49.545 49.76 49.618 ;
      RECT 47.868 49.499 49.806 49.572 ;
      RECT 47.914 49.453 49.852 49.526 ;
      RECT 47.96 49.407 49.898 49.48 ;
      RECT 48.006 49.361 49.944 49.434 ;
      RECT 48.052 49.315 49.99 49.388 ;
      RECT 48.098 49.269 50.036 49.342 ;
      RECT 48.144 49.223 50.082 49.296 ;
      RECT 48.19 49.177 50.128 49.25 ;
      RECT 48.236 49.131 50.174 49.204 ;
      RECT 48.282 49.085 50.22 49.158 ;
      RECT 48.328 49.039 50.266 49.112 ;
      RECT 48.374 48.993 50.312 49.066 ;
      RECT 48.42 48.947 50.358 49.02 ;
      RECT 48.466 48.901 50.404 48.974 ;
      RECT 48.512 48.855 50.45 48.928 ;
      RECT 48.558 48.809 50.496 48.882 ;
      RECT 48.604 48.763 50.542 48.836 ;
      RECT 48.65 48.717 50.588 48.79 ;
      RECT 48.696 48.671 50.634 48.744 ;
      RECT 48.742 48.625 50.68 48.698 ;
      RECT 48.788 48.579 50.726 48.652 ;
      RECT 48.834 48.533 50.772 48.606 ;
      RECT 48.88 48.487 50.818 48.56 ;
      RECT 48.926 48.441 50.864 48.514 ;
      RECT 48.972 48.395 50.91 48.468 ;
      RECT 49.018 48.349 50.956 48.422 ;
      RECT 49.064 48.303 51.002 48.376 ;
      RECT 49.11 48.257 51.048 48.33 ;
      RECT 49.156 48.211 51.094 48.284 ;
      RECT 49.202 48.165 51.14 48.238 ;
      RECT 49.248 48.119 51.186 48.192 ;
      RECT 49.294 48.073 51.232 48.146 ;
      RECT 49.34 48.027 51.278 48.1 ;
      RECT 49.386 47.981 51.324 48.054 ;
      RECT 49.432 47.935 51.37 48.008 ;
      RECT 49.478 47.889 51.416 47.962 ;
      RECT 49.524 47.843 51.462 47.916 ;
      RECT 49.57 47.797 51.508 47.87 ;
      RECT 49.616 47.751 51.554 47.824 ;
      RECT 49.662 47.705 51.6 47.778 ;
      RECT 49.708 47.659 51.646 47.732 ;
      RECT 49.754 47.613 51.692 47.686 ;
      RECT 49.8 47.567 51.738 47.64 ;
      RECT 49.846 47.521 51.784 47.594 ;
      RECT 49.892 47.475 51.83 47.548 ;
      RECT 49.938 47.429 51.876 47.502 ;
      RECT 49.984 47.383 51.922 47.456 ;
      RECT 50.03 47.337 51.968 47.41 ;
      RECT 50.076 47.291 52.014 47.364 ;
      RECT 50.122 47.245 52.06 47.318 ;
      RECT 50.168 47.199 52.106 47.272 ;
      RECT 50.214 47.153 52.152 47.226 ;
      RECT 50.26 47.107 52.198 47.18 ;
      RECT 50.306 47.061 52.244 47.134 ;
      RECT 50.352 47.015 52.29 47.088 ;
      RECT 50.398 46.969 52.336 47.042 ;
      RECT 50.444 46.923 52.382 46.996 ;
      RECT 50.49 46.877 52.428 46.95 ;
      RECT 50.536 46.831 52.474 46.904 ;
      RECT 50.582 46.785 52.52 46.858 ;
      RECT 50.628 46.739 52.566 46.812 ;
      RECT 50.674 46.693 52.612 46.766 ;
      RECT 50.72 46.647 52.658 46.72 ;
      RECT 50.766 46.601 52.704 46.674 ;
      RECT 50.812 46.555 52.75 46.628 ;
      RECT 50.858 46.509 52.796 46.582 ;
      RECT 50.904 46.463 52.842 46.536 ;
      RECT 50.95 46.417 52.888 46.49 ;
      RECT 50.996 46.371 52.934 46.444 ;
      RECT 51.042 46.325 52.98 46.398 ;
      RECT 51.088 46.279 53.026 46.352 ;
      RECT 51.134 46.233 53.072 46.306 ;
      RECT 51.18 46.187 53.118 46.26 ;
      RECT 51.226 46.141 53.164 46.214 ;
      RECT 51.272 46.095 53.21 46.168 ;
      RECT 51.318 46.049 53.256 46.122 ;
      RECT 51.364 46.003 53.302 46.076 ;
      RECT 51.41 45.957 53.348 46.03 ;
      RECT 51.456 45.911 53.394 45.984 ;
      RECT 51.502 45.865 53.44 45.938 ;
      RECT 51.548 45.819 53.486 45.892 ;
      RECT 51.594 45.773 53.532 45.846 ;
      RECT 51.64 45.727 53.578 45.8 ;
      RECT 51.686 45.681 53.624 45.754 ;
      RECT 51.732 45.635 53.67 45.708 ;
      RECT 51.778 45.589 53.716 45.662 ;
      RECT 51.824 45.543 53.762 45.616 ;
      RECT 51.87 45.497 53.808 45.57 ;
      RECT 51.916 45.451 53.854 45.524 ;
      RECT 51.962 45.405 53.9 45.478 ;
      RECT 52.008 45.359 53.946 45.432 ;
      RECT 52.054 45.313 53.992 45.386 ;
      RECT 52.1 45.267 54.038 45.34 ;
      RECT 52.146 45.221 54.084 45.294 ;
      RECT 52.192 45.175 54.13 45.248 ;
      RECT 52.238 45.129 54.176 45.202 ;
      RECT 52.284 45.083 54.222 45.156 ;
      RECT 52.33 45.037 54.268 45.11 ;
      RECT 52.376 44.991 54.314 45.064 ;
      RECT 52.422 44.945 54.36 45.018 ;
      RECT 52.468 44.899 54.406 44.972 ;
      RECT 52.514 44.853 54.452 44.926 ;
      RECT 52.56 44.807 54.498 44.88 ;
      RECT 52.606 44.761 54.544 44.834 ;
      RECT 52.652 44.715 54.59 44.788 ;
      RECT 52.698 44.669 54.636 44.742 ;
      RECT 52.744 44.623 54.682 44.696 ;
      RECT 52.79 44.577 54.728 44.65 ;
      RECT 52.836 44.531 54.774 44.604 ;
      RECT 52.882 44.485 54.82 44.558 ;
      RECT 52.928 44.439 54.866 44.512 ;
      RECT 52.974 44.393 54.912 44.466 ;
      RECT 53.02 44.347 54.958 44.42 ;
      RECT 53.066 44.301 55.004 44.374 ;
      RECT 53.112 44.255 55.05 44.328 ;
      RECT 53.158 44.209 55.096 44.282 ;
      RECT 53.204 44.163 55.142 44.236 ;
      RECT 53.25 44.117 55.188 44.19 ;
      RECT 53.296 44.071 55.234 44.144 ;
      RECT 53.342 44.025 55.28 44.098 ;
      RECT 53.388 43.979 55.326 44.052 ;
      RECT 53.434 43.933 55.372 44.006 ;
      RECT 53.48 43.887 55.418 43.96 ;
      RECT 53.526 43.841 55.464 43.914 ;
      RECT 53.572 43.795 55.51 43.868 ;
      RECT 53.618 43.749 55.556 43.822 ;
      RECT 53.664 43.703 55.602 43.776 ;
      RECT 53.71 43.657 55.648 43.73 ;
      RECT 53.756 43.611 55.694 43.684 ;
      RECT 53.802 43.565 55.74 43.638 ;
      RECT 53.848 43.519 55.786 43.592 ;
      RECT 53.894 43.473 55.832 43.546 ;
      RECT 53.94 43.427 55.878 43.5 ;
      RECT 53.986 43.381 55.924 43.454 ;
      RECT 54.032 43.335 55.97 43.408 ;
      RECT 54.078 43.289 56.016 43.362 ;
      RECT 54.124 43.243 56.062 43.316 ;
      RECT 54.17 43.197 56.108 43.27 ;
      RECT 54.216 43.151 56.154 43.224 ;
      RECT 54.262 43.105 56.2 43.178 ;
      RECT 54.308 43.059 56.246 43.132 ;
      RECT 54.354 43.013 56.292 43.086 ;
      RECT 54.4 42.967 56.338 43.04 ;
      RECT 54.446 42.921 56.384 42.994 ;
      RECT 54.492 42.875 56.43 42.948 ;
      RECT 54.538 42.829 56.476 42.902 ;
      RECT 54.584 42.783 56.522 42.856 ;
      RECT 54.63 42.737 56.568 42.81 ;
      RECT 54.676 42.691 56.614 42.764 ;
      RECT 54.722 42.645 56.66 42.718 ;
      RECT 54.768 42.599 56.706 42.672 ;
      RECT 54.814 42.553 56.752 42.626 ;
      RECT 54.86 42.507 56.798 42.58 ;
      RECT 54.906 42.461 56.844 42.534 ;
      RECT 54.952 42.415 56.89 42.488 ;
      RECT 54.998 42.369 56.936 42.442 ;
      RECT 55.044 42.323 56.982 42.396 ;
      RECT 55.09 42.277 57.028 42.35 ;
      RECT 55.136 42.231 57.074 42.304 ;
      RECT 55.182 42.185 57.12 42.258 ;
      RECT 55.228 42.139 57.166 42.212 ;
      RECT 55.274 42.093 57.212 42.166 ;
      RECT 55.32 42.047 57.258 42.12 ;
      RECT 55.366 42.001 57.304 42.074 ;
      RECT 55.412 41.955 57.35 42.028 ;
      RECT 55.458 41.909 57.396 41.982 ;
      RECT 55.504 41.863 57.442 41.936 ;
      RECT 55.55 41.817 57.488 41.89 ;
      RECT 55.596 41.771 57.534 41.844 ;
      RECT 55.642 41.725 57.58 41.798 ;
      RECT 55.688 41.679 57.626 41.752 ;
      RECT 55.734 41.633 57.672 41.706 ;
      RECT 55.78 41.587 57.718 41.66 ;
      RECT 55.826 41.541 57.764 41.614 ;
      RECT 55.872 41.495 57.81 41.568 ;
      RECT 55.918 41.449 57.856 41.522 ;
      RECT 55.964 41.403 57.902 41.476 ;
      RECT 56.01 41.357 57.948 41.43 ;
      RECT 56.056 41.311 57.994 41.384 ;
      RECT 56.102 41.265 58.04 41.338 ;
      RECT 56.148 41.219 58.086 41.292 ;
      RECT 56.194 41.173 58.132 41.246 ;
      RECT 56.24 41.127 58.178 41.2 ;
      RECT 56.286 41.081 58.224 41.154 ;
      RECT 56.332 41.035 58.27 41.108 ;
      RECT 56.378 40.989 58.316 41.062 ;
      RECT 56.424 40.943 58.362 41.016 ;
      RECT 56.47 40.897 58.408 40.97 ;
      RECT 56.516 40.851 58.454 40.924 ;
      RECT 56.562 40.805 58.5 40.878 ;
      RECT 56.608 40.759 58.546 40.832 ;
      RECT 56.654 40.713 58.592 40.786 ;
      RECT 56.7 40.667 58.638 40.74 ;
      RECT 56.746 40.621 58.684 40.694 ;
      RECT 56.792 40.575 58.73 40.648 ;
      RECT 56.838 40.529 58.776 40.602 ;
      RECT 56.884 40.483 58.822 40.556 ;
      RECT 56.93 40.437 58.868 40.51 ;
      RECT 56.976 40.391 58.914 40.464 ;
      RECT 57.022 40.345 58.96 40.418 ;
      RECT 57.068 40.299 59.006 40.372 ;
      RECT 57.114 40.253 59.052 40.326 ;
      RECT 57.16 40.207 59.098 40.28 ;
      RECT 57.206 40.161 59.144 40.234 ;
      RECT 57.252 40.115 59.19 40.188 ;
      RECT 57.298 40.069 59.236 40.142 ;
      RECT 57.344 40.023 59.282 40.096 ;
      RECT 57.39 39.977 59.328 40.05 ;
      RECT 57.436 39.931 59.374 40.004 ;
      RECT 57.482 39.885 59.42 39.958 ;
      RECT 57.528 39.839 59.466 39.912 ;
      RECT 57.574 39.793 59.512 39.866 ;
      RECT 57.62 39.747 59.558 39.82 ;
      RECT 57.666 39.701 59.604 39.774 ;
      RECT 57.712 39.655 59.65 39.728 ;
      RECT 57.758 39.609 59.696 39.682 ;
      RECT 57.804 39.563 59.742 39.636 ;
      RECT 57.85 39.517 59.788 39.59 ;
      RECT 57.896 39.471 59.834 39.544 ;
      RECT 57.942 39.425 59.88 39.498 ;
      RECT 57.988 39.379 59.926 39.452 ;
      RECT 58.034 39.333 59.972 39.406 ;
      RECT 58.08 39.287 60.018 39.36 ;
      RECT 58.126 39.241 60.064 39.314 ;
      RECT 58.172 39.195 60.11 39.268 ;
      RECT 58.218 39.149 60.156 39.222 ;
      RECT 58.264 39.103 60.202 39.176 ;
      RECT 58.31 39.057 60.248 39.13 ;
      RECT 58.356 39.011 60.294 39.084 ;
      RECT 58.402 38.965 60.34 39.038 ;
      RECT 58.448 38.919 60.386 38.992 ;
      RECT 58.494 38.873 60.432 38.946 ;
      RECT 58.54 38.827 60.478 38.9 ;
      RECT 58.586 38.781 60.524 38.854 ;
      RECT 58.632 38.735 60.57 38.808 ;
      RECT 58.678 38.689 60.616 38.762 ;
      RECT 58.724 38.643 60.662 38.716 ;
      RECT 58.77 38.597 60.708 38.67 ;
      RECT 58.816 38.551 60.754 38.624 ;
      RECT 58.862 38.505 60.8 38.578 ;
      RECT 58.908 38.459 60.846 38.532 ;
      RECT 58.954 38.413 60.892 38.486 ;
      RECT 59 38.367 60.938 38.44 ;
      RECT 59.046 38.321 60.984 38.394 ;
      RECT 59.092 38.275 61.03 38.348 ;
      RECT 59.138 38.229 61.076 38.302 ;
      RECT 59.184 38.183 61.122 38.256 ;
      RECT 59.23 38.137 61.168 38.21 ;
      RECT 59.276 38.091 61.214 38.164 ;
      RECT 59.322 38.045 61.26 38.118 ;
      RECT 59.368 37.999 61.306 38.072 ;
      RECT 59.414 37.953 61.352 38.026 ;
      RECT 59.46 37.907 61.398 37.98 ;
      RECT 59.506 37.861 61.444 37.934 ;
      RECT 59.552 37.815 61.49 37.888 ;
      RECT 59.598 37.769 61.536 37.842 ;
      RECT 59.644 37.723 61.582 37.796 ;
      RECT 59.69 37.677 61.628 37.75 ;
      RECT 59.736 37.631 61.674 37.704 ;
      RECT 59.782 37.585 61.72 37.658 ;
      RECT 59.828 37.539 61.766 37.612 ;
      RECT 59.874 37.493 61.812 37.566 ;
      RECT 59.92 37.447 61.858 37.52 ;
      RECT 59.966 37.401 61.904 37.474 ;
      RECT 60.012 37.355 61.95 37.428 ;
      RECT 60.058 37.309 61.996 37.382 ;
      RECT 60.104 37.263 62.042 37.336 ;
      RECT 60.15 37.217 62.088 37.29 ;
      RECT 60.196 37.171 62.134 37.244 ;
      RECT 60.242 37.125 62.18 37.198 ;
      RECT 60.288 37.079 62.226 37.152 ;
      RECT 60.334 37.033 62.272 37.106 ;
      RECT 60.38 36.987 62.318 37.06 ;
      RECT 60.426 36.941 62.364 37.014 ;
      RECT 60.472 36.895 62.41 36.968 ;
      RECT 60.518 36.849 62.456 36.922 ;
      RECT 60.564 36.803 62.502 36.876 ;
      RECT 60.61 36.757 62.548 36.83 ;
      RECT 60.656 36.711 62.594 36.784 ;
      RECT 60.702 36.665 62.64 36.738 ;
      RECT 60.748 36.619 62.686 36.692 ;
      RECT 60.794 36.573 62.732 36.646 ;
      RECT 60.84 36.527 62.778 36.6 ;
      RECT 60.886 36.481 62.824 36.554 ;
      RECT 60.932 36.435 62.87 36.508 ;
      RECT 60.978 36.389 62.916 36.462 ;
      RECT 61.024 36.343 62.962 36.416 ;
      RECT 61.07 36.297 63.008 36.37 ;
      RECT 61.116 36.251 63.054 36.324 ;
      RECT 61.162 36.205 63.1 36.278 ;
      RECT 63.094 34.296 63.1 36.278 ;
      RECT 61.208 36.159 63.146 36.232 ;
      RECT 63.095 34.272 63.146 36.232 ;
      RECT 61.254 36.113 63.192 36.186 ;
      RECT 63.141 34.226 63.192 36.186 ;
      RECT 61.3 36.067 63.238 36.14 ;
      RECT 63.187 34.18 63.238 36.14 ;
      RECT 61.346 36.021 63.284 36.094 ;
      RECT 63.233 34.134 63.284 36.094 ;
      RECT 61.392 35.975 63.33 36.048 ;
      RECT 63.279 34.088 63.33 36.048 ;
      RECT 61.438 35.929 63.376 36.002 ;
      RECT 63.325 34.042 63.376 36.002 ;
      RECT 61.484 35.883 63.422 35.956 ;
      RECT 63.371 33.996 63.422 35.956 ;
      RECT 61.53 35.837 63.468 35.91 ;
      RECT 63.417 33.95 63.468 35.91 ;
      RECT 61.576 35.791 63.514 35.864 ;
      RECT 63.463 33.904 63.514 35.864 ;
      RECT 61.622 35.745 63.56 35.818 ;
      RECT 63.509 33.858 63.56 35.818 ;
      RECT 61.668 35.699 63.606 35.772 ;
      RECT 63.555 33.812 63.606 35.772 ;
      RECT 61.714 35.653 63.652 35.726 ;
      RECT 63.601 33.766 63.652 35.726 ;
      RECT 61.76 35.607 63.698 35.68 ;
      RECT 63.647 33.72 63.698 35.68 ;
      RECT 61.806 35.561 63.744 35.634 ;
      RECT 63.693 33.674 63.744 35.634 ;
      RECT 61.852 35.515 63.79 35.588 ;
      RECT 63.739 33.628 63.79 35.588 ;
      RECT 61.898 35.469 63.836 35.542 ;
      RECT 63.785 33.582 63.836 35.542 ;
      RECT 61.944 35.423 63.882 35.496 ;
      RECT 63.831 33.536 63.882 35.496 ;
      RECT 61.99 35.377 63.928 35.45 ;
      RECT 63.877 33.49 63.928 35.45 ;
      RECT 62.036 35.331 63.974 35.404 ;
      RECT 63.923 33.444 63.974 35.404 ;
      RECT 62.082 35.285 64.02 35.358 ;
      RECT 63.969 33.398 64.02 35.358 ;
      RECT 62.128 35.239 64.066 35.312 ;
      RECT 64.015 33.352 64.066 35.312 ;
      RECT 62.174 35.193 64.112 35.266 ;
      RECT 64.061 33.306 64.112 35.266 ;
      RECT 62.22 35.147 64.158 35.22 ;
      RECT 64.107 33.26 64.158 35.22 ;
      RECT 62.266 35.101 64.204 35.174 ;
      RECT 64.153 33.214 64.204 35.174 ;
      RECT 62.312 35.055 64.25 35.128 ;
      RECT 64.199 33.168 64.25 35.128 ;
      RECT 62.358 35.009 64.296 35.082 ;
      RECT 64.245 33.122 64.296 35.082 ;
      RECT 62.404 34.963 64.342 35.036 ;
      RECT 64.291 33.076 64.342 35.036 ;
      RECT 62.45 34.917 64.388 34.99 ;
      RECT 64.337 33.03 64.388 34.99 ;
      RECT 62.496 34.871 64.434 34.944 ;
      RECT 64.383 32.984 64.434 34.944 ;
      RECT 62.542 34.825 64.48 34.898 ;
      RECT 64.429 32.938 64.48 34.898 ;
      RECT 62.588 34.779 64.526 34.852 ;
      RECT 64.475 32.892 64.526 34.852 ;
      RECT 62.634 34.733 64.572 34.806 ;
      RECT 64.521 32.846 64.572 34.806 ;
      RECT 62.68 34.687 64.618 34.76 ;
      RECT 64.567 32.8 64.618 34.76 ;
      RECT 62.726 34.641 64.664 34.714 ;
      RECT 64.613 32.754 64.664 34.714 ;
      RECT 62.772 34.595 64.71 34.668 ;
      RECT 64.659 32.708 64.71 34.668 ;
      RECT 62.818 34.549 64.756 34.622 ;
      RECT 64.705 32.662 64.756 34.622 ;
      RECT 62.864 34.503 64.802 34.576 ;
      RECT 64.751 32.616 64.802 34.576 ;
      RECT 62.91 34.457 64.848 34.53 ;
      RECT 64.797 32.57 64.848 34.53 ;
      RECT 62.956 34.411 64.894 34.484 ;
      RECT 64.843 32.524 64.894 34.484 ;
      RECT 63.002 34.365 64.94 34.438 ;
      RECT 64.889 32.478 64.94 34.438 ;
      RECT 63.048 34.319 64.986 34.392 ;
      RECT 64.935 32.432 64.986 34.392 ;
      RECT 64.981 32.386 65.032 34.346 ;
      RECT 65.027 32.34 65.078 34.3 ;
      RECT 65.073 32.294 65.124 34.254 ;
      RECT 65.119 32.248 65.17 34.208 ;
      RECT 65.165 32.202 65.216 34.162 ;
      RECT 65.211 32.156 65.262 34.116 ;
      RECT 65.257 32.11 65.308 34.07 ;
      RECT 65.303 32.064 65.354 34.024 ;
      RECT 65.349 32.018 65.4 33.978 ;
      RECT 65.395 31.972 65.446 33.932 ;
      RECT 65.441 31.926 65.492 33.886 ;
      RECT 65.487 31.88 65.538 33.84 ;
      RECT 65.533 31.834 65.584 33.794 ;
      RECT 65.579 31.788 65.63 33.748 ;
      RECT 65.625 31.742 65.676 33.702 ;
      RECT 65.671 31.696 65.722 33.656 ;
      RECT 65.717 31.65 65.768 33.61 ;
      RECT 65.763 31.604 65.814 33.564 ;
      RECT 65.809 31.558 65.86 33.518 ;
      RECT 65.855 31.512 65.906 33.472 ;
      RECT 65.901 31.466 65.952 33.426 ;
      RECT 65.947 31.42 65.998 33.38 ;
      RECT 65.993 31.374 66.044 33.334 ;
      RECT 66.039 31.328 66.09 33.288 ;
      RECT 66.085 31.282 66.136 33.242 ;
      RECT 66.131 31.236 66.182 33.196 ;
      RECT 66.177 31.19 66.228 33.15 ;
      RECT 66.223 31.144 66.274 33.104 ;
      RECT 66.269 31.098 66.32 33.058 ;
      RECT 66.315 31.052 66.366 33.012 ;
      RECT 66.361 31.006 66.412 32.966 ;
      RECT 66.407 30.96 66.458 32.92 ;
      RECT 66.453 30.914 66.504 32.874 ;
      RECT 66.499 30.868 66.55 32.828 ;
      RECT 66.545 30.822 66.596 32.782 ;
      RECT 66.591 30.776 66.642 32.736 ;
      RECT 66.637 30.73 66.688 32.69 ;
      RECT 66.683 30.684 66.734 32.644 ;
      RECT 66.729 30.638 66.78 32.598 ;
      RECT 66.775 30.592 66.826 32.552 ;
      RECT 66.821 30.546 66.872 32.506 ;
      RECT 66.867 30.5 66.918 32.46 ;
      RECT 66.913 30.454 66.964 32.414 ;
      RECT 66.959 30.408 67.01 32.368 ;
      RECT 67.005 30.362 67.056 32.322 ;
      RECT 67.051 30.316 67.102 32.276 ;
      RECT 67.097 30.27 67.148 32.23 ;
      RECT 67.143 30.224 67.194 32.184 ;
      RECT 67.189 30.178 67.24 32.138 ;
      RECT 67.235 30.132 67.286 32.092 ;
      RECT 67.281 30.086 67.332 32.046 ;
      RECT 67.327 30.04 67.378 32 ;
      RECT 67.373 29.994 67.424 31.954 ;
      RECT 67.419 29.948 67.47 31.908 ;
      RECT 67.465 29.902 67.516 31.862 ;
      RECT 67.511 29.856 67.562 31.816 ;
      RECT 67.557 29.81 67.608 31.77 ;
      RECT 67.603 29.764 67.654 31.724 ;
      RECT 67.649 29.718 67.7 31.678 ;
      RECT 67.695 29.672 67.746 31.632 ;
      RECT 67.741 29.626 67.792 31.586 ;
      RECT 67.787 29.58 67.838 31.54 ;
      RECT 67.833 29.534 67.884 31.494 ;
      RECT 67.879 29.488 67.93 31.448 ;
      RECT 67.925 29.442 67.976 31.402 ;
      RECT 67.971 29.396 68.022 31.356 ;
      RECT 68.017 29.352 68.068 31.31 ;
      RECT 68.06 29.33 68.114 31.264 ;
      RECT 68.06 29.33 68.16 31.218 ;
      RECT 68.06 29.33 68.206 31.172 ;
      RECT 68.06 29.33 68.252 31.126 ;
      RECT 68.06 29.33 68.298 31.08 ;
      RECT 68.06 29.33 68.344 31.034 ;
      RECT 68.06 29.33 68.39 30.988 ;
      RECT 68.06 29.33 68.436 30.942 ;
      RECT 68.06 29.33 68.482 30.896 ;
      RECT 68.06 29.33 68.528 30.85 ;
      RECT 68.06 29.33 68.574 30.804 ;
      RECT 68.06 29.33 68.62 30.758 ;
      RECT 68.06 29.33 68.666 30.712 ;
      RECT 68.06 29.33 68.712 30.666 ;
      RECT 68.06 29.33 68.758 30.62 ;
      RECT 68.06 29.33 68.804 30.574 ;
      RECT 68.06 29.33 68.85 30.528 ;
      RECT 68.06 29.33 68.896 30.482 ;
      RECT 68.06 29.33 68.942 30.436 ;
      RECT 68.06 29.33 68.988 30.39 ;
      RECT 68.06 29.33 69.034 30.344 ;
      RECT 68.06 29.33 69.08 30.298 ;
      RECT 68.06 29.33 69.126 30.252 ;
      RECT 68.06 29.33 69.172 30.206 ;
      RECT 67.235 30.132 69.185 30.176 ;
      RECT 68.06 29.33 110 30.17 ;
      RECT 42.83 74.787 43.67 110 ;
      RECT 42.83 74.787 43.716 75.912 ;
      RECT 42.83 74.787 43.762 75.866 ;
      RECT 42.83 74.787 43.808 75.82 ;
      RECT 42.83 74.787 43.854 75.774 ;
      RECT 42.83 74.787 43.9 75.728 ;
      RECT 42.83 74.787 43.946 75.682 ;
      RECT 42.83 74.787 43.992 75.636 ;
      RECT 42.83 74.787 44.038 75.59 ;
      RECT 42.83 74.787 44.084 75.544 ;
      RECT 42.83 74.787 44.13 75.498 ;
      RECT 42.83 74.787 44.176 75.452 ;
      RECT 42.83 74.787 44.222 75.406 ;
      RECT 42.83 74.787 44.268 75.36 ;
      RECT 42.83 74.787 44.314 75.314 ;
      RECT 42.83 74.787 44.36 75.268 ;
      RECT 42.83 74.787 44.406 75.222 ;
      RECT 42.83 74.787 44.452 75.176 ;
      RECT 42.83 74.787 44.498 75.13 ;
      RECT 42.83 74.787 44.544 75.084 ;
      RECT 42.83 74.787 44.59 75.038 ;
      RECT 42.83 74.787 44.636 74.992 ;
      RECT 42.83 74.787 44.682 74.946 ;
      RECT 42.83 74.787 44.728 74.9 ;
      RECT 42.83 74.787 44.774 74.854 ;
      RECT 42.876 74.741 44.82 74.808 ;
      RECT 44.762 72.855 44.82 74.808 ;
      RECT 42.922 74.695 44.866 74.762 ;
      RECT 44.808 72.809 44.866 74.762 ;
      RECT 42.968 74.649 44.912 74.716 ;
      RECT 44.854 72.763 44.912 74.716 ;
      RECT 43.014 74.603 44.958 74.67 ;
      RECT 44.9 72.717 44.958 74.67 ;
      RECT 43.06 74.557 45.004 74.624 ;
      RECT 44.946 72.671 45.004 74.624 ;
      RECT 43.106 74.511 45.05 74.578 ;
      RECT 44.992 72.625 45.05 74.578 ;
      RECT 43.152 74.465 45.096 74.532 ;
      RECT 45.038 72.579 45.096 74.532 ;
      RECT 43.198 74.419 45.142 74.486 ;
      RECT 45.084 72.533 45.142 74.486 ;
      RECT 43.244 74.373 45.188 74.44 ;
      RECT 45.13 72.487 45.188 74.44 ;
      RECT 43.29 74.327 45.234 74.394 ;
      RECT 45.176 72.441 45.234 74.394 ;
      RECT 43.336 74.281 45.28 74.348 ;
      RECT 45.222 72.395 45.28 74.348 ;
      RECT 43.382 74.235 45.326 74.302 ;
      RECT 45.268 72.349 45.326 74.302 ;
      RECT 43.428 74.189 45.372 74.256 ;
      RECT 45.314 72.303 45.372 74.256 ;
      RECT 43.474 74.143 45.418 74.21 ;
      RECT 45.36 72.257 45.418 74.21 ;
      RECT 43.52 74.097 45.464 74.164 ;
      RECT 45.406 72.211 45.464 74.164 ;
      RECT 43.566 74.051 45.51 74.118 ;
      RECT 45.452 72.165 45.51 74.118 ;
      RECT 43.612 74.005 45.556 74.072 ;
      RECT 45.498 72.119 45.556 74.072 ;
      RECT 43.658 73.959 45.602 74.026 ;
      RECT 45.544 72.073 45.602 74.026 ;
      RECT 43.704 73.913 45.648 73.98 ;
      RECT 45.59 72.027 45.648 73.98 ;
      RECT 43.75 73.867 45.694 73.934 ;
      RECT 45.636 71.981 45.694 73.934 ;
      RECT 43.796 73.821 45.74 73.888 ;
      RECT 45.682 71.935 45.74 73.888 ;
      RECT 43.842 73.775 45.786 73.842 ;
      RECT 45.728 71.889 45.786 73.842 ;
      RECT 43.888 73.729 45.832 73.796 ;
      RECT 45.774 71.843 45.832 73.796 ;
      RECT 43.934 73.683 45.878 73.75 ;
      RECT 45.82 71.797 45.878 73.75 ;
      RECT 43.98 73.637 45.924 73.704 ;
      RECT 45.866 71.751 45.924 73.704 ;
      RECT 44.026 73.591 45.97 73.658 ;
      RECT 45.912 71.705 45.97 73.658 ;
      RECT 44.072 73.545 46.016 73.612 ;
      RECT 45.958 71.659 46.016 73.612 ;
      RECT 44.118 73.499 46.062 73.566 ;
      RECT 46.004 71.613 46.062 73.566 ;
      RECT 44.164 73.453 46.108 73.52 ;
      RECT 46.05 71.567 46.108 73.52 ;
      RECT 44.21 73.407 46.154 73.474 ;
      RECT 46.096 71.521 46.154 73.474 ;
      RECT 44.256 73.361 46.2 73.428 ;
      RECT 46.142 71.475 46.2 73.428 ;
      RECT 44.302 73.315 46.246 73.382 ;
      RECT 46.188 71.429 46.246 73.382 ;
      RECT 44.348 73.269 46.292 73.336 ;
      RECT 46.234 71.383 46.292 73.336 ;
      RECT 44.394 73.223 46.338 73.29 ;
      RECT 46.28 71.337 46.338 73.29 ;
      RECT 44.44 73.177 46.384 73.244 ;
      RECT 46.326 71.291 46.384 73.244 ;
      RECT 44.486 73.131 46.43 73.198 ;
      RECT 46.372 71.245 46.43 73.198 ;
      RECT 44.532 73.085 46.476 73.152 ;
      RECT 46.418 71.199 46.476 73.152 ;
      RECT 44.578 73.039 46.522 73.106 ;
      RECT 46.464 71.153 46.522 73.106 ;
      RECT 44.624 72.993 46.568 73.06 ;
      RECT 46.51 71.107 46.568 73.06 ;
      RECT 44.67 72.947 46.614 73.014 ;
      RECT 46.556 71.061 46.614 73.014 ;
      RECT 44.716 72.901 46.66 72.968 ;
      RECT 46.602 71.015 46.66 72.968 ;
      RECT 46.648 70.969 46.706 72.922 ;
      RECT 46.694 70.923 46.752 72.876 ;
      RECT 46.74 70.877 46.798 72.83 ;
      RECT 46.786 70.831 46.844 72.784 ;
      RECT 46.832 70.785 46.89 72.738 ;
      RECT 46.878 70.739 46.936 72.692 ;
      RECT 46.924 70.693 46.982 72.646 ;
      RECT 46.97 70.647 47.028 72.6 ;
      RECT 47.016 70.601 47.074 72.554 ;
      RECT 47.062 70.555 47.12 72.508 ;
      RECT 47.108 70.509 47.166 72.462 ;
      RECT 47.154 70.463 47.212 72.416 ;
      RECT 47.2 70.417 47.258 72.37 ;
      RECT 47.246 70.371 47.304 72.324 ;
      RECT 47.292 70.325 47.35 72.278 ;
      RECT 47.338 70.279 47.396 72.232 ;
      RECT 47.384 70.233 47.442 72.186 ;
      RECT 47.43 70.187 47.488 72.14 ;
      RECT 47.476 70.141 47.534 72.094 ;
      RECT 47.522 70.095 47.58 72.048 ;
      RECT 47.568 70.049 47.626 72.002 ;
      RECT 47.614 70.003 47.672 71.956 ;
      RECT 47.66 69.957 47.718 71.91 ;
      RECT 47.706 69.911 47.764 71.864 ;
      RECT 47.752 69.865 47.81 71.818 ;
      RECT 47.798 69.819 47.856 71.772 ;
      RECT 47.844 69.773 47.902 71.726 ;
      RECT 47.89 69.727 47.948 71.68 ;
      RECT 47.936 69.681 47.994 71.634 ;
      RECT 47.982 69.635 48.04 71.588 ;
      RECT 48.028 69.589 48.086 71.542 ;
      RECT 48.074 69.543 48.132 71.496 ;
      RECT 48.12 69.497 48.178 71.45 ;
      RECT 48.166 69.451 48.224 71.404 ;
      RECT 48.212 69.405 48.27 71.358 ;
      RECT 48.258 69.359 48.316 71.312 ;
      RECT 48.304 69.313 48.362 71.266 ;
      RECT 48.35 69.267 48.408 71.22 ;
      RECT 48.396 69.221 48.454 71.174 ;
      RECT 48.442 69.175 48.5 71.128 ;
      RECT 48.488 69.129 48.546 71.082 ;
      RECT 48.534 69.083 48.592 71.036 ;
      RECT 48.58 69.037 48.638 70.99 ;
      RECT 48.626 68.991 48.684 70.944 ;
      RECT 48.672 68.945 48.73 70.898 ;
      RECT 48.718 68.899 48.776 70.852 ;
      RECT 48.764 68.853 48.822 70.806 ;
      RECT 48.81 68.807 48.868 70.76 ;
      RECT 48.856 68.761 48.914 70.714 ;
      RECT 48.902 68.715 48.96 70.668 ;
      RECT 48.948 68.669 49.006 70.622 ;
      RECT 48.994 68.623 49.052 70.576 ;
      RECT 49.04 68.577 49.098 70.53 ;
      RECT 49.086 68.531 49.144 70.484 ;
      RECT 49.132 68.485 49.19 70.438 ;
      RECT 49.178 68.439 49.236 70.392 ;
      RECT 49.224 68.393 49.282 70.346 ;
      RECT 49.27 68.347 49.328 70.3 ;
      RECT 49.316 68.301 49.374 70.254 ;
      RECT 49.362 68.255 49.42 70.208 ;
      RECT 49.408 68.209 49.466 70.162 ;
      RECT 49.454 68.163 49.512 70.116 ;
      RECT 49.5 68.117 49.558 70.07 ;
      RECT 49.546 68.071 49.604 70.024 ;
      RECT 49.592 68.025 49.65 69.978 ;
      RECT 49.638 67.979 49.696 69.932 ;
      RECT 49.684 67.933 49.742 69.886 ;
      RECT 49.73 67.887 49.788 69.84 ;
      RECT 49.776 67.841 49.834 69.794 ;
      RECT 49.822 67.795 49.88 69.748 ;
      RECT 49.868 67.749 49.926 69.702 ;
      RECT 49.914 67.703 49.972 69.656 ;
      RECT 49.96 67.657 50.018 69.61 ;
      RECT 50.006 67.611 50.064 69.564 ;
      RECT 50.052 67.565 50.11 69.518 ;
      RECT 50.098 67.519 50.156 69.472 ;
      RECT 50.144 67.473 50.202 69.426 ;
      RECT 50.19 67.427 50.248 69.38 ;
      RECT 50.236 67.381 50.294 69.334 ;
      RECT 50.282 67.335 50.34 69.288 ;
      RECT 50.328 67.289 50.386 69.242 ;
      RECT 50.374 67.243 50.432 69.196 ;
      RECT 50.42 67.197 50.478 69.15 ;
      RECT 50.466 67.151 50.524 69.104 ;
      RECT 50.512 67.105 50.57 69.058 ;
      RECT 50.558 67.059 50.616 69.012 ;
      RECT 50.604 67.013 50.662 68.966 ;
      RECT 50.65 66.967 50.708 68.92 ;
      RECT 50.696 66.921 50.754 68.874 ;
      RECT 50.742 66.875 50.8 68.828 ;
      RECT 50.788 66.829 50.846 68.782 ;
      RECT 50.834 66.783 50.892 68.736 ;
      RECT 50.88 66.737 50.938 68.69 ;
      RECT 50.926 66.691 50.984 68.644 ;
      RECT 50.972 66.645 51.03 68.598 ;
      RECT 51.018 66.599 51.076 68.552 ;
      RECT 51.064 66.553 51.122 68.506 ;
      RECT 51.11 66.507 51.168 68.46 ;
      RECT 51.156 66.461 51.214 68.414 ;
      RECT 51.202 66.415 51.26 68.368 ;
      RECT 51.248 66.369 51.306 68.322 ;
      RECT 51.294 66.323 51.352 68.276 ;
      RECT 51.34 66.277 51.398 68.23 ;
      RECT 51.386 66.231 51.444 68.184 ;
      RECT 51.432 66.185 51.49 68.138 ;
      RECT 51.478 66.139 51.536 68.092 ;
      RECT 51.524 66.093 51.582 68.046 ;
      RECT 51.57 66.047 51.628 68 ;
      RECT 51.616 66.001 51.674 67.954 ;
      RECT 51.662 65.955 51.72 67.908 ;
      RECT 51.708 65.909 51.766 67.862 ;
      RECT 51.754 65.863 51.812 67.816 ;
      RECT 51.8 65.817 51.858 67.77 ;
      RECT 51.846 65.771 51.904 67.724 ;
      RECT 51.892 65.725 51.95 67.678 ;
      RECT 51.938 65.679 51.996 67.632 ;
      RECT 51.984 65.633 52.042 67.586 ;
      RECT 52.03 65.587 52.088 67.54 ;
      RECT 52.076 65.541 52.134 67.494 ;
      RECT 52.122 65.495 52.18 67.448 ;
      RECT 52.168 65.449 52.226 67.402 ;
      RECT 52.214 65.403 52.272 67.356 ;
      RECT 52.26 65.357 52.318 67.31 ;
      RECT 52.306 65.311 52.364 67.264 ;
      RECT 52.352 65.265 52.41 67.218 ;
      RECT 52.398 65.219 52.456 67.172 ;
      RECT 52.444 65.173 52.502 67.126 ;
      RECT 52.49 65.127 52.548 67.08 ;
      RECT 52.536 65.081 52.594 67.034 ;
      RECT 52.582 65.035 52.64 66.988 ;
      RECT 52.628 64.989 52.686 66.942 ;
      RECT 52.674 64.943 52.732 66.896 ;
      RECT 52.72 64.897 52.778 66.85 ;
      RECT 52.766 64.851 52.824 66.804 ;
      RECT 52.812 64.805 52.87 66.758 ;
      RECT 52.858 64.759 52.916 66.712 ;
      RECT 52.904 64.713 52.962 66.666 ;
      RECT 52.95 64.667 53.008 66.62 ;
      RECT 52.996 64.621 53.054 66.574 ;
      RECT 53.042 64.575 53.1 66.528 ;
      RECT 53.088 64.529 53.146 66.482 ;
      RECT 53.134 64.483 53.192 66.436 ;
      RECT 53.18 64.437 53.238 66.39 ;
      RECT 53.226 64.391 53.284 66.344 ;
      RECT 53.272 64.345 53.33 66.298 ;
      RECT 53.318 64.299 53.376 66.252 ;
      RECT 53.364 64.253 53.422 66.206 ;
      RECT 53.41 64.207 53.468 66.16 ;
      RECT 53.456 64.161 53.514 66.114 ;
      RECT 53.502 64.115 53.56 66.068 ;
      RECT 53.548 64.069 53.606 66.022 ;
      RECT 53.594 64.023 53.652 65.976 ;
      RECT 53.64 63.977 53.698 65.93 ;
      RECT 53.686 63.931 53.744 65.884 ;
      RECT 53.732 63.885 53.79 65.838 ;
      RECT 53.778 63.839 53.836 65.792 ;
      RECT 53.824 63.793 53.882 65.746 ;
      RECT 53.87 63.747 53.928 65.7 ;
      RECT 53.916 63.701 53.974 65.654 ;
      RECT 53.962 63.655 54.02 65.608 ;
      RECT 54.008 63.609 54.066 65.562 ;
      RECT 54.054 63.563 54.112 65.516 ;
      RECT 54.1 63.517 54.158 65.47 ;
      RECT 54.146 63.471 54.204 65.424 ;
      RECT 54.192 63.425 54.25 65.378 ;
      RECT 54.238 63.379 54.296 65.332 ;
      RECT 54.284 63.333 54.342 65.286 ;
      RECT 54.33 63.287 54.388 65.24 ;
      RECT 54.376 63.241 54.434 65.194 ;
      RECT 54.422 63.195 54.48 65.148 ;
      RECT 54.468 63.149 54.526 65.102 ;
      RECT 54.514 63.103 54.572 65.056 ;
      RECT 54.56 63.057 54.618 65.01 ;
      RECT 54.606 63.011 54.664 64.964 ;
      RECT 54.652 62.965 54.71 64.918 ;
      RECT 54.698 62.919 54.756 64.872 ;
      RECT 54.744 62.873 54.802 64.826 ;
      RECT 54.79 62.827 54.848 64.78 ;
      RECT 54.836 62.781 54.894 64.734 ;
      RECT 54.882 62.735 54.94 64.688 ;
      RECT 54.928 62.689 54.986 64.642 ;
      RECT 54.974 62.643 55.032 64.596 ;
      RECT 55.02 62.597 55.078 64.55 ;
      RECT 55.066 62.551 55.124 64.504 ;
      RECT 55.112 62.505 55.17 64.458 ;
      RECT 55.158 62.459 55.216 64.412 ;
      RECT 55.204 62.413 55.262 64.366 ;
      RECT 55.25 62.367 55.308 64.32 ;
      RECT 55.296 62.321 55.354 64.274 ;
      RECT 55.342 62.275 55.4 64.228 ;
      RECT 55.388 62.229 55.446 64.182 ;
      RECT 55.434 62.183 55.492 64.136 ;
      RECT 55.48 62.137 55.538 64.09 ;
      RECT 55.526 62.091 55.584 64.044 ;
      RECT 55.572 62.045 55.63 63.998 ;
      RECT 55.618 61.999 55.67 63.955 ;
      RECT 55.664 61.953 55.716 63.912 ;
      RECT 55.71 61.907 55.762 63.866 ;
      RECT 55.756 61.861 55.808 63.82 ;
      RECT 55.802 61.815 55.854 63.774 ;
      RECT 55.848 61.769 55.9 63.728 ;
      RECT 55.894 61.723 55.946 63.682 ;
      RECT 55.94 61.677 55.992 63.636 ;
      RECT 55.986 61.631 56.038 63.59 ;
      RECT 56.032 61.585 56.084 63.544 ;
      RECT 56.078 61.539 56.13 63.498 ;
      RECT 56.124 61.493 56.176 63.452 ;
      RECT 56.17 61.447 56.222 63.406 ;
      RECT 56.216 61.401 56.268 63.36 ;
      RECT 56.262 61.355 56.314 63.314 ;
      RECT 56.308 61.309 56.36 63.268 ;
      RECT 56.354 61.263 56.406 63.222 ;
      RECT 56.4 61.217 56.452 63.176 ;
      RECT 56.446 61.171 56.498 63.13 ;
      RECT 56.492 61.125 56.544 63.084 ;
      RECT 56.538 61.079 56.59 63.038 ;
      RECT 56.584 61.033 56.636 62.992 ;
      RECT 56.63 60.987 56.682 62.946 ;
      RECT 56.676 60.941 56.728 62.9 ;
      RECT 56.722 60.895 56.774 62.854 ;
      RECT 56.768 60.849 56.82 62.808 ;
      RECT 56.814 60.803 56.866 62.762 ;
      RECT 56.86 60.757 56.912 62.716 ;
      RECT 56.906 60.711 56.958 62.67 ;
      RECT 56.952 60.665 57.004 62.624 ;
      RECT 56.998 60.619 57.05 62.578 ;
      RECT 57.044 60.573 57.096 62.532 ;
      RECT 57.09 60.527 57.142 62.486 ;
      RECT 57.136 60.481 57.188 62.44 ;
      RECT 57.182 60.435 57.234 62.394 ;
      RECT 57.228 60.389 57.28 62.348 ;
      RECT 57.274 60.343 57.326 62.302 ;
      RECT 57.32 60.297 57.372 62.256 ;
      RECT 57.366 60.251 57.418 62.21 ;
      RECT 57.412 60.205 57.464 62.164 ;
      RECT 57.458 60.159 57.51 62.118 ;
      RECT 57.504 60.113 57.556 62.072 ;
      RECT 57.55 60.067 57.602 62.026 ;
      RECT 57.596 60.021 57.648 61.98 ;
      RECT 57.642 59.975 57.694 61.934 ;
      RECT 57.688 59.929 57.74 61.888 ;
      RECT 57.734 59.883 57.786 61.842 ;
      RECT 57.78 59.837 57.832 61.796 ;
      RECT 57.826 59.791 57.878 61.75 ;
      RECT 57.872 59.745 57.924 61.704 ;
      RECT 57.918 59.699 57.97 61.658 ;
      RECT 57.964 59.653 58.016 61.612 ;
      RECT 58.01 59.607 58.062 61.566 ;
      RECT 58.056 59.561 58.108 61.52 ;
      RECT 58.102 59.515 58.154 61.474 ;
      RECT 58.148 59.469 58.2 61.428 ;
      RECT 58.194 59.423 58.246 61.382 ;
      RECT 58.24 59.377 58.292 61.336 ;
      RECT 58.286 59.331 58.338 61.29 ;
      RECT 58.332 59.285 58.384 61.244 ;
      RECT 58.378 59.239 58.43 61.198 ;
      RECT 58.424 59.193 58.476 61.152 ;
      RECT 58.47 59.147 58.522 61.106 ;
      RECT 58.516 59.101 58.568 61.06 ;
      RECT 58.562 59.055 58.614 61.014 ;
      RECT 58.608 59.009 58.66 60.968 ;
      RECT 58.654 58.963 58.706 60.922 ;
      RECT 58.7 58.917 58.752 60.876 ;
      RECT 58.746 58.871 58.798 60.83 ;
      RECT 58.792 58.825 58.844 60.784 ;
      RECT 58.838 58.779 58.89 60.738 ;
      RECT 58.884 58.733 58.936 60.692 ;
      RECT 58.93 58.687 58.982 60.646 ;
      RECT 58.976 58.641 59.028 60.6 ;
      RECT 59.022 58.595 59.074 60.554 ;
      RECT 59.068 58.549 59.12 60.508 ;
      RECT 59.114 58.503 59.166 60.462 ;
      RECT 59.16 58.457 59.212 60.416 ;
      RECT 59.206 58.411 59.258 60.37 ;
      RECT 59.252 58.365 59.304 60.324 ;
      RECT 59.298 58.319 59.35 60.278 ;
      RECT 59.344 58.273 59.396 60.232 ;
      RECT 59.39 58.227 59.442 60.186 ;
      RECT 59.436 58.181 59.488 60.14 ;
      RECT 59.482 58.135 59.534 60.094 ;
      RECT 59.528 58.089 59.58 60.048 ;
      RECT 59.574 58.043 59.626 60.002 ;
      RECT 59.62 57.997 59.672 59.956 ;
      RECT 59.666 57.951 59.718 59.91 ;
      RECT 59.712 57.905 59.764 59.864 ;
      RECT 59.758 57.859 59.81 59.818 ;
      RECT 59.804 57.813 59.856 59.772 ;
      RECT 59.85 57.767 59.902 59.726 ;
      RECT 59.896 57.721 59.948 59.68 ;
      RECT 59.942 57.675 59.994 59.634 ;
      RECT 59.988 57.629 60.04 59.588 ;
      RECT 60.034 57.583 60.086 59.542 ;
      RECT 60.08 57.537 60.132 59.496 ;
      RECT 60.126 57.491 60.178 59.45 ;
      RECT 60.172 57.445 60.224 59.404 ;
      RECT 60.218 57.399 60.27 59.358 ;
      RECT 60.264 57.353 60.316 59.312 ;
      RECT 60.31 57.307 60.362 59.266 ;
      RECT 60.356 57.261 60.408 59.22 ;
      RECT 60.402 57.215 60.454 59.174 ;
      RECT 60.448 57.169 60.5 59.128 ;
      RECT 60.494 57.123 60.546 59.082 ;
      RECT 60.54 57.077 60.592 59.036 ;
      RECT 60.586 57.031 60.638 58.99 ;
      RECT 60.632 56.985 60.684 58.944 ;
      RECT 60.678 56.939 60.73 58.898 ;
      RECT 60.724 56.893 60.776 58.852 ;
      RECT 60.77 56.847 60.822 58.806 ;
      RECT 60.816 56.801 60.868 58.76 ;
      RECT 60.862 56.755 60.914 58.714 ;
      RECT 60.908 56.709 60.96 58.668 ;
      RECT 60.954 56.663 61.006 58.622 ;
      RECT 61 56.617 61.052 58.576 ;
      RECT 61.046 56.571 61.098 58.53 ;
      RECT 61.092 56.525 61.144 58.484 ;
      RECT 61.138 56.479 61.19 58.438 ;
      RECT 61.184 56.433 61.236 58.392 ;
      RECT 61.23 56.387 61.282 58.346 ;
      RECT 61.276 56.341 61.328 58.3 ;
      RECT 61.322 56.295 61.374 58.254 ;
      RECT 61.368 56.249 61.42 58.208 ;
      RECT 61.414 56.203 61.466 58.162 ;
      RECT 61.46 56.157 61.512 58.116 ;
      RECT 61.506 56.111 61.558 58.07 ;
      RECT 61.552 56.065 61.604 58.024 ;
      RECT 61.598 56.019 61.65 57.978 ;
      RECT 61.644 55.973 61.696 57.932 ;
      RECT 61.69 55.927 61.742 57.886 ;
      RECT 61.736 55.881 61.788 57.84 ;
      RECT 61.782 55.835 61.834 57.794 ;
      RECT 61.828 55.789 61.88 57.748 ;
      RECT 61.874 55.743 61.926 57.702 ;
      RECT 61.92 55.697 61.972 57.656 ;
      RECT 61.966 55.651 62.018 57.61 ;
      RECT 62.012 55.605 62.064 57.564 ;
      RECT 62.058 55.559 62.11 57.518 ;
      RECT 62.104 55.513 62.156 57.472 ;
      RECT 62.15 55.467 62.202 57.426 ;
      RECT 62.196 55.421 62.248 57.38 ;
      RECT 62.242 55.375 62.294 57.334 ;
      RECT 62.288 55.329 62.34 57.288 ;
      RECT 62.334 55.283 62.386 57.242 ;
      RECT 62.38 55.237 62.432 57.196 ;
      RECT 62.426 55.191 62.478 57.15 ;
      RECT 62.472 55.145 62.524 57.104 ;
      RECT 62.518 55.099 62.57 57.058 ;
      RECT 62.564 55.053 62.616 57.012 ;
      RECT 62.61 55.007 62.662 56.966 ;
      RECT 62.656 54.961 62.708 56.92 ;
      RECT 62.702 54.915 62.754 56.874 ;
      RECT 62.748 54.869 62.8 56.828 ;
      RECT 62.794 54.823 62.846 56.782 ;
      RECT 62.84 54.777 62.892 56.736 ;
      RECT 62.886 54.731 62.938 56.69 ;
      RECT 62.932 54.685 62.984 56.644 ;
      RECT 62.978 54.639 63.03 56.598 ;
      RECT 63.024 54.593 63.076 56.552 ;
      RECT 63.07 54.547 63.122 56.506 ;
      RECT 63.116 54.501 63.168 56.46 ;
      RECT 63.162 54.455 63.214 56.414 ;
      RECT 63.208 54.409 63.26 56.368 ;
      RECT 63.254 54.363 63.306 56.322 ;
      RECT 63.3 54.317 63.352 56.276 ;
      RECT 63.346 54.271 63.398 56.23 ;
      RECT 63.392 54.225 63.444 56.184 ;
      RECT 63.438 54.179 63.49 56.138 ;
      RECT 63.484 54.133 63.536 56.092 ;
      RECT 63.53 54.087 63.582 56.046 ;
      RECT 63.576 54.041 63.628 56 ;
      RECT 63.622 53.995 63.674 55.954 ;
      RECT 63.668 53.949 63.72 55.908 ;
      RECT 63.714 53.903 63.766 55.862 ;
      RECT 63.76 53.857 63.812 55.816 ;
      RECT 63.806 53.811 63.858 55.77 ;
      RECT 63.852 53.765 63.904 55.724 ;
      RECT 63.898 53.719 63.95 55.678 ;
      RECT 63.944 53.673 63.996 55.632 ;
      RECT 63.99 53.627 64.042 55.586 ;
      RECT 64.036 53.581 64.088 55.54 ;
      RECT 64.082 53.535 64.134 55.494 ;
      RECT 64.128 53.489 64.18 55.448 ;
      RECT 64.174 53.443 64.226 55.402 ;
      RECT 64.22 53.397 64.272 55.356 ;
      RECT 64.266 53.351 64.318 55.31 ;
      RECT 64.312 53.305 64.364 55.264 ;
      RECT 64.358 53.259 64.41 55.218 ;
      RECT 64.404 53.213 64.456 55.172 ;
      RECT 64.45 53.167 64.502 55.126 ;
      RECT 64.496 53.121 64.548 55.08 ;
      RECT 64.542 53.075 64.594 55.034 ;
      RECT 64.588 53.029 64.64 54.988 ;
      RECT 64.634 52.983 64.686 54.942 ;
      RECT 64.68 52.937 64.732 54.896 ;
      RECT 64.726 52.891 64.778 54.85 ;
      RECT 64.772 52.845 64.824 54.804 ;
      RECT 64.818 52.799 64.87 54.758 ;
      RECT 64.864 52.753 64.916 54.712 ;
      RECT 64.91 52.707 64.962 54.666 ;
      RECT 64.956 52.661 65.008 54.62 ;
      RECT 65.002 52.615 65.054 54.574 ;
      RECT 65.048 52.569 65.1 54.528 ;
      RECT 65.094 52.523 65.146 54.482 ;
      RECT 65.14 52.477 65.192 54.436 ;
      RECT 65.186 52.431 65.238 54.39 ;
      RECT 65.232 52.385 65.284 54.344 ;
      RECT 65.278 52.339 65.33 54.298 ;
      RECT 65.324 52.293 65.376 54.252 ;
      RECT 65.37 52.247 65.422 54.206 ;
      RECT 65.416 52.201 65.468 54.16 ;
      RECT 65.462 52.155 65.514 54.114 ;
      RECT 65.508 52.109 65.56 54.068 ;
      RECT 65.554 52.063 65.606 54.022 ;
      RECT 65.6 52.017 65.652 53.976 ;
      RECT 65.646 51.971 65.698 53.93 ;
      RECT 65.692 51.925 65.744 53.884 ;
      RECT 65.738 51.879 65.79 53.838 ;
      RECT 65.784 51.833 65.836 53.792 ;
      RECT 65.83 51.787 65.882 53.746 ;
      RECT 65.876 51.741 65.928 53.7 ;
      RECT 65.922 51.695 65.974 53.654 ;
      RECT 65.968 51.649 66.02 53.608 ;
      RECT 66.014 51.603 66.066 53.562 ;
      RECT 66.06 51.557 66.112 53.516 ;
      RECT 66.106 51.511 66.158 53.47 ;
      RECT 66.152 51.465 66.204 53.424 ;
      RECT 66.198 51.419 66.25 53.378 ;
      RECT 66.244 51.373 66.296 53.332 ;
      RECT 66.29 51.327 66.342 53.286 ;
      RECT 66.336 51.281 66.388 53.24 ;
      RECT 66.382 51.235 66.434 53.194 ;
      RECT 66.428 51.189 66.48 53.148 ;
      RECT 66.474 51.143 66.526 53.102 ;
      RECT 66.52 51.097 66.572 53.056 ;
      RECT 66.566 51.051 66.618 53.01 ;
      RECT 66.612 51.005 66.664 52.964 ;
      RECT 66.658 50.959 66.71 52.918 ;
      RECT 66.704 50.913 66.756 52.872 ;
      RECT 66.75 50.867 66.802 52.826 ;
      RECT 66.796 50.821 66.848 52.78 ;
      RECT 66.842 50.775 66.894 52.734 ;
      RECT 66.888 50.729 66.94 52.688 ;
      RECT 66.934 50.683 66.986 52.642 ;
      RECT 66.98 50.637 67.032 52.596 ;
      RECT 67.026 50.591 67.078 52.55 ;
      RECT 67.072 50.545 67.124 52.504 ;
      RECT 67.118 50.499 67.17 52.458 ;
      RECT 67.164 50.453 67.216 52.412 ;
      RECT 67.21 50.407 67.262 52.366 ;
      RECT 67.256 50.361 67.308 52.32 ;
      RECT 67.302 50.315 67.354 52.274 ;
      RECT 67.348 50.269 67.4 52.228 ;
      RECT 67.394 50.223 67.446 52.182 ;
      RECT 67.44 50.177 67.492 52.136 ;
      RECT 67.486 50.131 67.538 52.09 ;
      RECT 67.532 50.085 67.584 52.044 ;
      RECT 67.578 50.039 67.63 51.998 ;
      RECT 67.624 49.993 67.676 51.952 ;
      RECT 67.67 49.947 67.722 51.906 ;
      RECT 67.716 49.901 67.768 51.86 ;
      RECT 67.762 49.855 67.814 51.814 ;
      RECT 67.808 49.809 67.86 51.768 ;
      RECT 67.854 49.763 67.906 51.722 ;
      RECT 67.9 49.717 67.952 51.676 ;
      RECT 67.946 49.671 67.998 51.63 ;
      RECT 67.992 49.625 68.044 51.584 ;
      RECT 68.038 49.579 68.09 51.538 ;
      RECT 68.084 49.533 68.136 51.492 ;
      RECT 68.13 49.487 68.182 51.446 ;
      RECT 68.176 49.441 68.228 51.4 ;
      RECT 68.222 49.395 68.274 51.354 ;
      RECT 68.268 49.349 68.32 51.308 ;
      RECT 68.314 49.303 68.366 51.262 ;
      RECT 68.36 49.257 68.412 51.216 ;
      RECT 68.406 49.211 68.458 51.17 ;
      RECT 68.452 49.165 68.504 51.124 ;
      RECT 68.498 49.119 68.55 51.078 ;
      RECT 68.544 49.073 68.596 51.032 ;
      RECT 68.59 49.027 68.642 50.986 ;
      RECT 68.636 48.981 68.688 50.94 ;
      RECT 68.682 48.935 68.734 50.894 ;
      RECT 68.728 48.889 68.78 50.848 ;
      RECT 68.774 48.843 68.826 50.802 ;
      RECT 68.82 48.797 68.872 50.756 ;
      RECT 68.866 48.751 68.918 50.71 ;
      RECT 68.912 48.705 68.964 50.664 ;
      RECT 68.958 48.659 69.01 50.618 ;
      RECT 69.004 48.613 69.056 50.572 ;
      RECT 69.05 48.567 69.102 50.526 ;
      RECT 69.096 48.521 69.148 50.48 ;
      RECT 69.142 48.475 69.194 50.434 ;
      RECT 69.188 48.429 69.24 50.388 ;
      RECT 69.234 48.383 69.286 50.342 ;
      RECT 69.28 48.337 69.332 50.296 ;
      RECT 69.326 48.291 69.378 50.25 ;
      RECT 69.372 48.245 69.424 50.204 ;
      RECT 69.418 48.199 69.47 50.158 ;
      RECT 69.464 48.153 69.516 50.112 ;
      RECT 69.51 48.107 69.562 50.066 ;
      RECT 69.556 48.061 69.608 50.02 ;
      RECT 69.602 48.015 69.654 49.974 ;
      RECT 69.648 47.969 69.7 49.928 ;
      RECT 69.694 47.923 69.746 49.882 ;
      RECT 69.74 47.877 69.792 49.836 ;
      RECT 69.786 47.831 69.838 49.79 ;
      RECT 69.832 47.802 69.884 49.744 ;
      RECT 69.845 47.772 69.93 49.698 ;
      RECT 69.891 47.726 69.976 49.652 ;
      RECT 69.937 47.68 70.022 49.606 ;
      RECT 69.983 47.634 70.068 49.56 ;
      RECT 70.029 47.588 70.114 49.514 ;
      RECT 70.075 47.542 70.16 49.468 ;
      RECT 70.121 47.496 70.206 49.422 ;
      RECT 70.167 47.45 70.252 49.376 ;
      RECT 70.213 47.404 70.298 49.33 ;
      RECT 70.259 47.358 70.344 49.284 ;
      RECT 70.305 47.312 70.39 49.238 ;
      RECT 70.351 47.266 70.436 49.192 ;
      RECT 70.397 47.22 70.482 49.146 ;
      RECT 70.443 47.174 70.528 49.1 ;
      RECT 70.489 47.128 70.574 49.054 ;
      RECT 70.535 47.082 70.62 49.008 ;
      RECT 70.581 47.036 70.666 48.962 ;
      RECT 70.627 46.99 70.712 48.916 ;
      RECT 70.673 46.944 70.758 48.87 ;
      RECT 70.719 46.898 70.804 48.824 ;
      RECT 70.765 46.852 70.85 48.778 ;
      RECT 70.811 46.806 70.896 48.732 ;
      RECT 70.857 46.76 70.942 48.686 ;
      RECT 70.903 46.714 70.988 48.64 ;
      RECT 70.949 46.668 71.034 48.594 ;
      RECT 70.995 46.622 71.08 48.548 ;
      RECT 71.041 46.576 71.126 48.502 ;
      RECT 71.087 46.53 71.172 48.456 ;
      RECT 71.133 46.484 71.218 48.41 ;
      RECT 71.179 46.438 71.264 48.364 ;
      RECT 71.225 46.392 71.31 48.318 ;
      RECT 71.271 46.346 71.356 48.272 ;
      RECT 71.317 46.3 71.402 48.226 ;
      RECT 71.363 46.254 71.448 48.18 ;
      RECT 71.409 46.208 71.494 48.134 ;
      RECT 71.455 46.162 71.54 48.088 ;
      RECT 71.501 46.116 71.586 48.042 ;
      RECT 71.547 46.07 71.632 47.996 ;
      RECT 71.593 46.024 71.678 47.95 ;
      RECT 71.639 45.978 71.724 47.904 ;
      RECT 71.685 45.932 71.77 47.858 ;
      RECT 71.731 45.886 71.816 47.812 ;
      RECT 71.777 45.84 71.862 47.766 ;
      RECT 71.823 45.794 71.908 47.72 ;
      RECT 71.869 45.748 71.954 47.674 ;
      RECT 71.915 45.702 72 47.628 ;
      RECT 71.961 45.656 72.046 47.582 ;
      RECT 72.007 45.61 72.092 47.536 ;
      RECT 72.053 45.564 72.138 47.49 ;
      RECT 72.099 45.518 72.184 47.444 ;
      RECT 72.145 45.472 72.23 47.398 ;
      RECT 72.191 45.426 72.276 47.352 ;
      RECT 72.237 45.38 72.322 47.306 ;
      RECT 72.283 45.334 72.368 47.26 ;
      RECT 72.329 45.288 72.414 47.214 ;
      RECT 72.375 45.242 72.46 47.168 ;
      RECT 72.421 45.196 72.506 47.122 ;
      RECT 72.467 45.15 72.552 47.076 ;
      RECT 72.513 45.104 72.598 47.03 ;
      RECT 72.559 45.058 72.644 46.984 ;
      RECT 72.605 45.012 72.69 46.938 ;
      RECT 72.651 44.966 72.736 46.892 ;
      RECT 72.697 44.92 72.782 46.846 ;
      RECT 72.743 44.874 72.828 46.8 ;
      RECT 72.789 44.828 72.874 46.754 ;
      RECT 72.835 44.782 72.92 46.708 ;
      RECT 72.881 44.736 72.966 46.662 ;
      RECT 72.927 44.69 73.012 46.616 ;
      RECT 72.973 44.644 73.058 46.57 ;
      RECT 73.019 44.598 73.104 46.524 ;
      RECT 73.065 44.552 73.15 46.478 ;
      RECT 73.111 44.506 73.196 46.432 ;
      RECT 73.157 44.46 73.242 46.386 ;
      RECT 73.203 44.414 73.288 46.34 ;
      RECT 73.249 44.368 73.334 46.294 ;
      RECT 73.295 44.322 73.38 46.248 ;
      RECT 73.341 44.276 73.426 46.202 ;
      RECT 73.387 44.23 73.472 46.156 ;
      RECT 73.433 44.184 73.518 46.11 ;
      RECT 73.479 44.138 73.564 46.064 ;
      RECT 73.525 44.092 73.61 46.018 ;
      RECT 73.571 44.046 73.656 45.972 ;
      RECT 73.617 44 73.702 45.926 ;
      RECT 73.663 43.954 73.748 45.88 ;
      RECT 73.709 43.908 73.794 45.834 ;
      RECT 73.755 43.862 73.84 45.788 ;
      RECT 73.801 43.816 73.886 45.742 ;
      RECT 73.847 43.77 73.932 45.696 ;
      RECT 73.893 43.724 73.978 45.65 ;
      RECT 73.939 43.678 74.024 45.604 ;
      RECT 73.985 43.632 74.07 45.558 ;
      RECT 74.031 43.586 74.116 45.512 ;
      RECT 74.077 43.54 74.162 45.466 ;
      RECT 74.123 43.494 74.208 45.42 ;
      RECT 74.169 43.448 74.254 45.374 ;
      RECT 74.215 43.402 74.3 45.328 ;
      RECT 74.261 43.356 74.346 45.282 ;
      RECT 74.307 43.31 74.392 45.236 ;
      RECT 74.353 43.264 74.438 45.19 ;
      RECT 74.399 43.218 74.484 45.144 ;
      RECT 74.445 43.172 74.53 45.098 ;
      RECT 74.491 43.126 74.576 45.052 ;
      RECT 74.537 43.08 74.622 45.006 ;
      RECT 74.583 43.034 74.668 44.96 ;
      RECT 74.629 42.988 74.714 44.914 ;
      RECT 74.675 42.942 74.76 44.868 ;
      RECT 74.721 42.896 74.806 44.822 ;
      RECT 74.767 42.852 74.852 44.776 ;
      RECT 74.81 42.83 74.898 44.73 ;
      RECT 74.81 42.83 74.944 44.684 ;
      RECT 74.81 42.83 74.99 44.638 ;
      RECT 74.81 42.83 75.036 44.592 ;
      RECT 74.81 42.83 75.082 44.546 ;
      RECT 74.81 42.83 75.128 44.5 ;
      RECT 74.81 42.83 75.174 44.454 ;
      RECT 74.81 42.83 75.22 44.408 ;
      RECT 74.81 42.83 75.266 44.362 ;
      RECT 74.81 42.83 75.312 44.316 ;
      RECT 74.81 42.83 75.358 44.27 ;
      RECT 74.81 42.83 75.404 44.224 ;
      RECT 74.81 42.83 75.45 44.178 ;
      RECT 74.81 42.83 75.496 44.132 ;
      RECT 74.81 42.83 75.542 44.086 ;
      RECT 74.81 42.83 75.588 44.04 ;
      RECT 74.81 42.83 75.634 43.994 ;
      RECT 74.81 42.83 75.68 43.948 ;
      RECT 74.81 42.83 75.726 43.902 ;
      RECT 74.81 42.83 75.772 43.856 ;
      RECT 74.81 42.83 75.818 43.81 ;
      RECT 74.81 42.83 75.864 43.764 ;
      RECT 73.939 43.678 75.91 43.718 ;
      RECT 74.81 42.83 75.935 43.682 ;
      RECT 74.81 42.83 110 43.67 ;
      RECT 76.595 61.272 78.35 61.273 ;
      RECT 76.641 61.226 78.35 61.273 ;
      RECT 76.641 61.226 78.396 61.227 ;
      RECT 76.687 61.18 78.396 61.227 ;
      RECT 76.687 61.18 78.442 61.181 ;
      RECT 76.733 61.134 78.442 61.181 ;
      RECT 76.733 61.134 78.488 61.135 ;
      RECT 76.779 61.088 78.488 61.135 ;
      RECT 76.779 61.088 78.534 61.089 ;
      RECT 76.825 61.042 78.534 61.089 ;
      RECT 76.825 61.042 78.58 61.043 ;
      RECT 76.871 60.996 78.58 61.043 ;
      RECT 76.871 60.996 78.626 60.997 ;
      RECT 76.917 60.95 78.626 60.997 ;
      RECT 76.917 60.95 78.672 60.951 ;
      RECT 76.963 60.904 78.672 60.951 ;
      RECT 76.963 60.904 78.718 60.905 ;
      RECT 77.009 60.858 78.718 60.905 ;
      RECT 77.009 60.858 78.764 60.859 ;
      RECT 77.055 60.812 78.764 60.859 ;
      RECT 77.055 60.812 78.81 60.813 ;
      RECT 77.101 60.766 78.81 60.813 ;
      RECT 77.101 60.766 78.856 60.767 ;
      RECT 77.147 60.72 78.856 60.767 ;
      RECT 77.147 60.72 78.902 60.721 ;
      RECT 77.193 60.674 78.902 60.721 ;
      RECT 77.193 60.674 78.948 60.675 ;
      RECT 77.239 60.628 78.948 60.675 ;
      RECT 77.239 60.628 78.994 60.629 ;
      RECT 77.285 60.582 78.994 60.629 ;
      RECT 77.285 60.582 79.04 60.583 ;
      RECT 77.331 60.536 79.04 60.583 ;
      RECT 77.331 60.536 79.086 60.537 ;
      RECT 77.377 60.49 79.086 60.537 ;
      RECT 77.377 60.49 79.132 60.491 ;
      RECT 77.423 60.444 79.132 60.491 ;
      RECT 77.423 60.444 79.178 60.445 ;
      RECT 77.469 60.398 79.178 60.445 ;
      RECT 77.469 60.398 79.224 60.399 ;
      RECT 77.515 60.352 79.224 60.399 ;
      RECT 77.515 60.352 79.27 60.353 ;
      RECT 77.561 60.306 79.27 60.353 ;
      RECT 77.561 60.306 79.316 60.307 ;
      RECT 77.607 60.26 79.316 60.307 ;
      RECT 77.607 60.26 79.362 60.261 ;
      RECT 77.653 60.214 79.362 60.261 ;
      RECT 77.653 60.214 79.408 60.215 ;
      RECT 77.699 60.168 79.408 60.215 ;
      RECT 77.699 60.168 79.454 60.169 ;
      RECT 77.745 60.122 79.454 60.169 ;
      RECT 77.745 60.122 79.5 60.123 ;
      RECT 77.791 60.076 79.5 60.123 ;
      RECT 77.791 60.076 79.546 60.077 ;
      RECT 77.837 60.03 79.546 60.077 ;
      RECT 77.837 60.03 79.592 60.031 ;
      RECT 77.883 59.984 79.592 60.031 ;
      RECT 77.883 59.984 79.638 59.985 ;
      RECT 77.929 59.938 79.638 59.985 ;
      RECT 77.929 59.938 79.684 59.939 ;
      RECT 77.975 59.892 79.684 59.939 ;
      RECT 77.975 59.892 79.73 59.893 ;
      RECT 78.021 59.846 79.73 59.893 ;
      RECT 78.021 59.846 79.776 59.847 ;
      RECT 78.067 59.8 79.776 59.847 ;
      RECT 78.067 59.8 79.822 59.801 ;
      RECT 78.113 59.754 79.822 59.801 ;
      RECT 78.113 59.754 79.868 59.755 ;
      RECT 78.159 59.708 79.868 59.755 ;
      RECT 78.159 59.708 79.914 59.709 ;
      RECT 78.205 59.662 79.914 59.709 ;
      RECT 78.205 59.662 79.96 59.663 ;
      RECT 78.251 59.616 79.96 59.663 ;
      RECT 78.251 59.616 80.006 59.617 ;
      RECT 78.297 59.57 80.006 59.617 ;
      RECT 78.297 59.57 80.052 59.571 ;
      RECT 78.343 59.524 80.052 59.571 ;
      RECT 78.343 59.524 80.098 59.525 ;
      RECT 78.389 59.478 80.098 59.525 ;
      RECT 78.389 59.478 80.144 59.479 ;
      RECT 78.435 59.432 80.144 59.479 ;
      RECT 78.435 59.432 80.19 59.433 ;
      RECT 78.481 59.386 80.19 59.433 ;
      RECT 78.481 59.386 80.236 59.387 ;
      RECT 78.527 59.34 80.236 59.387 ;
      RECT 78.527 59.34 80.282 59.341 ;
      RECT 78.573 59.294 80.282 59.341 ;
      RECT 78.573 59.294 80.328 59.295 ;
      RECT 78.619 59.248 80.328 59.295 ;
      RECT 78.619 59.248 80.374 59.249 ;
      RECT 78.665 59.202 80.374 59.249 ;
      RECT 78.665 59.202 80.42 59.203 ;
      RECT 78.711 59.156 80.42 59.203 ;
      RECT 78.711 59.156 80.466 59.157 ;
      RECT 78.757 59.11 80.466 59.157 ;
      RECT 78.757 59.11 80.512 59.111 ;
      RECT 78.803 59.064 80.512 59.111 ;
      RECT 78.803 59.064 80.558 59.065 ;
      RECT 78.849 59.018 80.558 59.065 ;
      RECT 78.849 59.018 80.604 59.019 ;
      RECT 78.895 58.972 80.604 59.019 ;
      RECT 78.895 58.972 80.65 58.973 ;
      RECT 78.941 58.926 80.65 58.973 ;
      RECT 78.941 58.926 80.696 58.927 ;
      RECT 78.987 58.88 80.696 58.927 ;
      RECT 78.987 58.88 80.742 58.881 ;
      RECT 79.033 58.834 80.742 58.881 ;
      RECT 79.033 58.834 80.788 58.835 ;
      RECT 79.079 58.788 80.788 58.835 ;
      RECT 79.079 58.788 80.834 58.789 ;
      RECT 79.125 58.742 80.834 58.789 ;
      RECT 79.125 58.742 80.88 58.743 ;
      RECT 79.171 58.696 80.88 58.743 ;
      RECT 79.171 58.696 80.926 58.697 ;
      RECT 79.217 58.65 80.926 58.697 ;
      RECT 79.217 58.65 80.972 58.651 ;
      RECT 79.263 58.604 80.972 58.651 ;
      RECT 79.263 58.604 81.018 58.605 ;
      RECT 79.309 58.558 81.018 58.605 ;
      RECT 79.309 58.558 81.064 58.559 ;
      RECT 79.355 58.512 81.064 58.559 ;
      RECT 79.355 58.512 81.11 58.513 ;
      RECT 79.401 58.466 81.11 58.513 ;
      RECT 79.401 58.466 81.156 58.467 ;
      RECT 79.447 58.42 81.156 58.467 ;
      RECT 79.447 58.42 81.202 58.421 ;
      RECT 79.493 58.374 81.202 58.421 ;
      RECT 79.493 58.374 81.248 58.375 ;
      RECT 79.539 58.328 81.248 58.375 ;
      RECT 79.539 58.328 81.294 58.329 ;
      RECT 79.585 58.282 81.294 58.329 ;
      RECT 79.585 58.282 81.34 58.283 ;
      RECT 79.631 58.236 81.34 58.283 ;
      RECT 79.631 58.236 81.386 58.237 ;
      RECT 79.677 58.19 81.386 58.237 ;
      RECT 79.677 58.19 81.432 58.191 ;
      RECT 79.723 58.144 81.432 58.191 ;
      RECT 79.723 58.144 81.478 58.145 ;
      RECT 79.769 58.098 81.478 58.145 ;
      RECT 79.769 58.098 81.524 58.099 ;
      RECT 79.815 58.052 81.524 58.099 ;
      RECT 79.815 58.052 81.57 58.053 ;
      RECT 79.861 58.006 81.57 58.053 ;
      RECT 79.861 58.006 81.616 58.007 ;
      RECT 79.907 57.96 81.662 57.961 ;
      RECT 79.953 57.914 81.708 57.915 ;
      RECT 79.999 57.868 81.754 57.869 ;
      RECT 80.045 57.822 81.8 57.823 ;
      RECT 80.091 57.776 81.846 57.777 ;
      RECT 80.137 57.73 81.892 57.731 ;
      RECT 80.183 57.684 81.938 57.685 ;
      RECT 80.229 57.638 81.984 57.639 ;
      RECT 80.275 57.592 82.03 57.593 ;
      RECT 80.321 57.546 82.076 57.547 ;
      RECT 80.367 57.5 82.122 57.501 ;
      RECT 80.413 57.454 82.168 57.455 ;
      RECT 80.459 57.408 82.214 57.409 ;
      RECT 80.505 57.362 82.26 57.363 ;
      RECT 80.551 57.316 82.306 57.317 ;
      RECT 80.597 57.27 82.352 57.271 ;
      RECT 80.643 57.224 82.398 57.225 ;
      RECT 56.33 81.537 57.17 110 ;
      RECT 56.33 81.537 57.216 82.407 ;
      RECT 56.33 81.537 57.262 82.361 ;
      RECT 56.33 81.537 57.308 82.315 ;
      RECT 56.33 81.537 57.354 82.269 ;
      RECT 56.33 81.537 57.4 82.223 ;
      RECT 56.33 81.537 57.446 82.177 ;
      RECT 56.33 81.537 57.492 82.131 ;
      RECT 56.33 81.537 57.538 82.085 ;
      RECT 56.33 81.537 57.584 82.039 ;
      RECT 56.33 81.537 57.63 81.993 ;
      RECT 56.33 81.537 57.676 81.947 ;
      RECT 56.33 81.537 57.722 81.901 ;
      RECT 56.33 81.537 57.768 81.855 ;
      RECT 56.33 81.537 57.814 81.809 ;
      RECT 56.33 81.537 57.86 81.763 ;
      RECT 56.33 81.537 57.906 81.717 ;
      RECT 56.33 81.537 57.952 81.671 ;
      RECT 56.33 81.537 57.998 81.625 ;
      RECT 56.376 81.491 58.044 81.579 ;
      RECT 56.422 81.445 58.09 81.533 ;
      RECT 56.468 81.399 58.136 81.487 ;
      RECT 56.514 81.353 58.182 81.441 ;
      RECT 56.56 81.307 58.228 81.395 ;
      RECT 56.606 81.261 58.274 81.349 ;
      RECT 56.652 81.215 58.32 81.303 ;
      RECT 56.698 81.169 58.366 81.257 ;
      RECT 56.744 81.123 58.412 81.211 ;
      RECT 56.79 81.077 58.458 81.165 ;
      RECT 56.836 81.031 58.504 81.119 ;
      RECT 56.882 80.985 58.55 81.073 ;
      RECT 56.928 80.939 58.596 81.027 ;
      RECT 56.974 80.893 58.642 80.981 ;
      RECT 57.02 80.847 58.688 80.935 ;
      RECT 57.066 80.801 58.734 80.889 ;
      RECT 57.112 80.755 58.78 80.843 ;
      RECT 57.158 80.709 58.826 80.797 ;
      RECT 57.204 80.663 58.872 80.751 ;
      RECT 57.25 80.617 58.918 80.705 ;
      RECT 57.296 80.571 58.964 80.659 ;
      RECT 57.342 80.525 59.01 80.613 ;
      RECT 57.388 80.479 59.056 80.567 ;
      RECT 57.434 80.433 59.102 80.521 ;
      RECT 57.48 80.387 59.148 80.475 ;
      RECT 57.526 80.341 59.194 80.429 ;
      RECT 57.572 80.295 59.24 80.383 ;
      RECT 57.618 80.249 59.286 80.337 ;
      RECT 57.664 80.203 59.332 80.291 ;
      RECT 57.71 80.157 59.378 80.245 ;
      RECT 57.756 80.111 59.424 80.199 ;
      RECT 57.802 80.065 59.47 80.153 ;
      RECT 57.848 80.019 59.516 80.107 ;
      RECT 57.894 79.973 59.562 80.061 ;
      RECT 57.94 79.927 59.608 80.015 ;
      RECT 57.986 79.881 59.654 79.969 ;
      RECT 58.032 79.835 59.7 79.923 ;
      RECT 58.078 79.789 59.746 79.877 ;
      RECT 58.124 79.743 59.792 79.831 ;
      RECT 58.17 79.697 59.838 79.785 ;
      RECT 58.216 79.651 59.884 79.739 ;
      RECT 58.262 79.605 59.93 79.693 ;
      RECT 58.308 79.559 59.976 79.647 ;
      RECT 58.354 79.513 60.022 79.601 ;
      RECT 58.4 79.467 60.068 79.555 ;
      RECT 58.446 79.421 60.114 79.509 ;
      RECT 58.492 79.375 60.16 79.463 ;
      RECT 58.538 79.329 60.206 79.417 ;
      RECT 58.584 79.283 60.252 79.371 ;
      RECT 58.63 79.237 60.298 79.325 ;
      RECT 58.676 79.191 60.344 79.279 ;
      RECT 58.722 79.145 60.39 79.233 ;
      RECT 58.768 79.099 60.436 79.187 ;
      RECT 58.814 79.053 60.482 79.141 ;
      RECT 58.86 79.007 60.528 79.095 ;
      RECT 58.906 78.961 60.574 79.049 ;
      RECT 58.952 78.915 60.62 79.003 ;
      RECT 58.998 78.869 60.666 78.957 ;
      RECT 59.044 78.823 60.712 78.911 ;
      RECT 59.09 78.777 60.758 78.865 ;
      RECT 59.136 78.731 60.804 78.819 ;
      RECT 59.182 78.685 60.85 78.773 ;
      RECT 59.228 78.639 60.896 78.727 ;
      RECT 59.274 78.593 60.942 78.681 ;
      RECT 59.32 78.547 60.988 78.635 ;
      RECT 59.366 78.501 61.034 78.589 ;
      RECT 59.412 78.455 61.08 78.543 ;
      RECT 59.458 78.409 61.126 78.497 ;
      RECT 59.504 78.363 61.172 78.451 ;
      RECT 59.55 78.317 61.218 78.405 ;
      RECT 59.596 78.271 61.264 78.359 ;
      RECT 59.642 78.225 61.31 78.313 ;
      RECT 59.688 78.179 61.356 78.267 ;
      RECT 59.734 78.133 61.402 78.221 ;
      RECT 59.78 78.087 61.448 78.175 ;
      RECT 59.826 78.041 61.494 78.129 ;
      RECT 59.872 77.995 61.54 78.083 ;
      RECT 59.918 77.949 61.586 78.037 ;
      RECT 59.964 77.903 61.632 77.991 ;
      RECT 60.01 77.857 61.678 77.945 ;
      RECT 60.056 77.811 61.724 77.899 ;
      RECT 60.102 77.765 61.77 77.853 ;
      RECT 60.148 77.719 61.816 77.807 ;
      RECT 60.194 77.673 61.862 77.761 ;
      RECT 60.24 77.627 61.908 77.715 ;
      RECT 60.286 77.581 61.954 77.669 ;
      RECT 60.332 77.535 62 77.623 ;
      RECT 60.378 77.489 62.046 77.577 ;
      RECT 60.424 77.443 62.092 77.531 ;
      RECT 60.47 77.397 62.138 77.485 ;
      RECT 60.516 77.351 62.184 77.439 ;
      RECT 60.562 77.305 62.23 77.393 ;
      RECT 60.608 77.259 62.276 77.347 ;
      RECT 60.654 77.213 62.322 77.301 ;
      RECT 60.7 77.167 62.368 77.255 ;
      RECT 60.746 77.121 62.414 77.209 ;
      RECT 60.792 77.075 62.46 77.163 ;
      RECT 60.838 77.029 62.506 77.117 ;
      RECT 60.884 76.983 62.552 77.071 ;
      RECT 60.93 76.937 62.598 77.025 ;
      RECT 60.976 76.891 62.644 76.979 ;
      RECT 61.022 76.845 62.69 76.933 ;
      RECT 61.068 76.799 62.736 76.887 ;
      RECT 61.114 76.753 62.782 76.841 ;
      RECT 61.16 76.707 62.828 76.795 ;
      RECT 61.206 76.661 62.874 76.749 ;
      RECT 61.252 76.615 62.92 76.703 ;
      RECT 61.298 76.569 62.966 76.657 ;
      RECT 61.344 76.523 63.012 76.611 ;
      RECT 61.39 76.477 63.058 76.565 ;
      RECT 61.436 76.431 63.104 76.519 ;
      RECT 61.436 76.431 63.15 76.473 ;
      RECT 61.482 76.385 63.17 76.44 ;
      RECT 61.528 76.339 63.216 76.407 ;
      RECT 61.574 76.293 63.262 76.361 ;
      RECT 61.62 76.247 63.308 76.315 ;
      RECT 61.666 76.201 63.354 76.269 ;
      RECT 61.712 76.155 63.4 76.223 ;
      RECT 61.758 76.109 63.446 76.177 ;
      RECT 61.804 76.063 63.492 76.131 ;
      RECT 61.85 76.017 63.538 76.085 ;
      RECT 61.896 75.971 63.584 76.039 ;
      RECT 61.942 75.925 63.63 75.993 ;
      RECT 61.988 75.879 63.676 75.947 ;
      RECT 62.034 75.833 63.722 75.901 ;
      RECT 62.08 75.787 63.768 75.855 ;
      RECT 62.126 75.741 63.814 75.809 ;
      RECT 62.172 75.695 63.86 75.763 ;
      RECT 62.218 75.649 63.906 75.717 ;
      RECT 62.264 75.603 63.952 75.671 ;
      RECT 62.31 75.557 63.998 75.625 ;
      RECT 62.356 75.511 64.044 75.579 ;
      RECT 62.402 75.465 64.09 75.533 ;
      RECT 62.448 75.419 64.136 75.487 ;
      RECT 62.494 75.373 64.182 75.441 ;
      RECT 62.54 75.327 64.228 75.395 ;
      RECT 62.586 75.281 64.274 75.349 ;
      RECT 62.632 75.235 64.32 75.303 ;
      RECT 62.678 75.189 64.366 75.257 ;
      RECT 62.724 75.143 64.412 75.211 ;
      RECT 62.77 75.097 64.458 75.165 ;
      RECT 62.816 75.051 64.504 75.119 ;
      RECT 62.862 75.005 64.55 75.073 ;
      RECT 62.908 74.959 64.596 75.027 ;
      RECT 62.954 74.913 64.642 74.981 ;
      RECT 63 74.867 64.688 74.935 ;
      RECT 63.046 74.821 64.734 74.889 ;
      RECT 63.092 74.775 64.78 74.843 ;
      RECT 63.138 74.729 64.826 74.797 ;
      RECT 63.184 74.683 64.872 74.751 ;
      RECT 63.23 74.637 64.918 74.705 ;
      RECT 63.276 74.591 64.964 74.659 ;
      RECT 63.322 74.545 65.01 74.613 ;
      RECT 63.368 74.499 65.056 74.567 ;
      RECT 63.414 74.453 65.102 74.521 ;
      RECT 63.46 74.407 65.148 74.475 ;
      RECT 63.506 74.361 65.194 74.429 ;
      RECT 63.552 74.315 65.24 74.383 ;
      RECT 63.598 74.269 65.286 74.337 ;
      RECT 63.644 74.223 65.332 74.291 ;
      RECT 63.69 74.177 65.378 74.245 ;
      RECT 63.736 74.131 65.424 74.199 ;
      RECT 63.782 74.085 65.47 74.153 ;
      RECT 63.828 74.039 65.516 74.107 ;
      RECT 63.874 73.993 65.562 74.061 ;
      RECT 63.92 73.947 65.608 74.015 ;
      RECT 63.966 73.901 65.654 73.969 ;
      RECT 64.012 73.855 65.7 73.923 ;
      RECT 64.058 73.809 65.746 73.877 ;
      RECT 64.104 73.763 65.792 73.831 ;
      RECT 64.15 73.717 65.838 73.785 ;
      RECT 64.196 73.671 65.884 73.739 ;
      RECT 64.242 73.625 65.93 73.693 ;
      RECT 64.288 73.579 65.976 73.647 ;
      RECT 64.334 73.533 66.022 73.601 ;
      RECT 64.38 73.487 66.068 73.555 ;
      RECT 64.426 73.441 66.114 73.509 ;
      RECT 64.472 73.395 66.16 73.463 ;
      RECT 64.518 73.349 66.206 73.417 ;
      RECT 64.564 73.303 66.252 73.371 ;
      RECT 64.61 73.257 66.298 73.325 ;
      RECT 64.656 73.211 66.344 73.279 ;
      RECT 64.702 73.165 66.39 73.233 ;
      RECT 64.748 73.119 66.436 73.187 ;
      RECT 64.794 73.073 66.482 73.141 ;
      RECT 64.84 73.027 66.528 73.095 ;
      RECT 64.886 72.981 66.574 73.049 ;
      RECT 64.932 72.935 66.62 73.003 ;
      RECT 64.978 72.889 66.666 72.957 ;
      RECT 65.024 72.843 66.712 72.911 ;
      RECT 65.07 72.797 66.758 72.865 ;
      RECT 65.116 72.751 66.804 72.819 ;
      RECT 65.162 72.705 66.85 72.773 ;
      RECT 65.208 72.659 66.896 72.727 ;
      RECT 65.254 72.613 66.942 72.681 ;
      RECT 65.3 72.567 66.988 72.635 ;
      RECT 65.346 72.521 67.034 72.589 ;
      RECT 65.392 72.475 67.08 72.543 ;
      RECT 65.438 72.429 67.126 72.497 ;
      RECT 65.484 72.383 67.172 72.451 ;
      RECT 65.53 72.337 67.218 72.405 ;
      RECT 65.576 72.291 67.264 72.359 ;
      RECT 65.622 72.245 67.31 72.313 ;
      RECT 65.668 72.199 67.356 72.267 ;
      RECT 65.714 72.153 67.402 72.221 ;
      RECT 65.76 72.107 67.448 72.175 ;
      RECT 65.806 72.061 67.494 72.129 ;
      RECT 65.852 72.015 67.54 72.083 ;
      RECT 65.898 71.969 67.586 72.037 ;
      RECT 65.944 71.923 67.632 71.991 ;
      RECT 65.99 71.877 67.678 71.945 ;
      RECT 66.036 71.831 67.724 71.899 ;
      RECT 66.082 71.785 67.77 71.853 ;
      RECT 66.128 71.739 67.816 71.807 ;
      RECT 66.174 71.693 67.862 71.761 ;
      RECT 66.22 71.647 67.908 71.715 ;
      RECT 66.266 71.601 67.954 71.669 ;
      RECT 66.312 71.555 68 71.623 ;
      RECT 66.358 71.509 68.046 71.577 ;
      RECT 66.404 71.463 68.092 71.531 ;
      RECT 66.45 71.417 68.138 71.485 ;
      RECT 66.496 71.371 68.184 71.439 ;
      RECT 66.542 71.325 68.23 71.393 ;
      RECT 66.588 71.279 68.276 71.347 ;
      RECT 66.634 71.233 68.322 71.301 ;
      RECT 66.68 71.187 68.368 71.255 ;
      RECT 66.726 71.141 68.414 71.209 ;
      RECT 66.772 71.095 68.46 71.163 ;
      RECT 66.818 71.049 68.506 71.117 ;
      RECT 66.864 71.003 68.552 71.071 ;
      RECT 66.91 70.957 68.598 71.025 ;
      RECT 66.956 70.911 68.644 70.979 ;
      RECT 67.002 70.865 68.69 70.933 ;
      RECT 67.048 70.819 68.736 70.887 ;
      RECT 67.094 70.773 68.782 70.841 ;
      RECT 67.14 70.727 68.828 70.795 ;
      RECT 67.186 70.681 68.874 70.749 ;
      RECT 67.232 70.635 68.92 70.703 ;
      RECT 67.278 70.589 68.966 70.657 ;
      RECT 67.324 70.543 69.012 70.611 ;
      RECT 67.37 70.497 69.058 70.565 ;
      RECT 67.416 70.451 69.104 70.519 ;
      RECT 67.462 70.405 69.15 70.473 ;
      RECT 67.508 70.359 69.196 70.427 ;
      RECT 67.554 70.313 69.242 70.381 ;
      RECT 67.6 70.267 69.288 70.335 ;
      RECT 67.646 70.221 69.334 70.289 ;
      RECT 67.692 70.175 69.38 70.243 ;
      RECT 67.738 70.129 69.426 70.197 ;
      RECT 67.784 70.083 69.472 70.151 ;
      RECT 67.83 70.037 69.518 70.105 ;
      RECT 67.876 69.991 69.564 70.059 ;
      RECT 67.922 69.945 69.61 70.013 ;
      RECT 67.968 69.899 69.656 69.967 ;
      RECT 68.014 69.853 69.702 69.921 ;
      RECT 68.06 69.807 69.748 69.875 ;
      RECT 68.106 69.761 69.794 69.829 ;
      RECT 68.152 69.715 69.84 69.783 ;
      RECT 68.198 69.669 69.886 69.737 ;
      RECT 68.244 69.623 69.932 69.691 ;
      RECT 68.29 69.577 69.978 69.645 ;
      RECT 68.336 69.531 70.024 69.599 ;
      RECT 68.382 69.485 70.07 69.553 ;
      RECT 68.428 69.439 70.116 69.507 ;
      RECT 68.474 69.393 70.162 69.461 ;
      RECT 68.52 69.347 70.208 69.415 ;
      RECT 68.566 69.301 70.254 69.369 ;
      RECT 68.612 69.255 70.3 69.323 ;
      RECT 68.658 69.209 70.346 69.277 ;
      RECT 68.704 69.163 70.392 69.231 ;
      RECT 68.75 69.117 70.438 69.185 ;
      RECT 68.796 69.071 70.484 69.139 ;
      RECT 68.842 69.025 70.53 69.093 ;
      RECT 68.888 68.979 70.576 69.047 ;
      RECT 68.934 68.933 70.622 69.001 ;
      RECT 68.98 68.887 70.668 68.955 ;
      RECT 69.026 68.841 70.714 68.909 ;
      RECT 69.072 68.795 70.76 68.863 ;
      RECT 69.118 68.749 70.806 68.817 ;
      RECT 69.164 68.703 70.852 68.771 ;
      RECT 69.21 68.657 70.898 68.725 ;
      RECT 69.256 68.611 70.944 68.679 ;
      RECT 69.302 68.565 70.99 68.633 ;
      RECT 69.348 68.519 71.036 68.587 ;
      RECT 69.394 68.473 71.082 68.541 ;
      RECT 69.44 68.427 71.128 68.495 ;
      RECT 69.486 68.381 71.174 68.449 ;
      RECT 69.532 68.335 71.22 68.403 ;
      RECT 69.578 68.289 71.266 68.357 ;
      RECT 69.624 68.243 71.312 68.311 ;
      RECT 69.67 68.197 71.358 68.265 ;
      RECT 69.716 68.151 71.404 68.219 ;
      RECT 69.762 68.105 71.45 68.173 ;
      RECT 69.808 68.059 71.496 68.127 ;
      RECT 69.854 68.013 71.542 68.081 ;
      RECT 69.9 67.967 71.588 68.035 ;
      RECT 69.946 67.921 71.634 67.989 ;
      RECT 69.992 67.875 71.68 67.943 ;
      RECT 70.038 67.829 71.726 67.897 ;
      RECT 70.084 67.783 71.772 67.851 ;
      RECT 70.13 67.737 71.818 67.805 ;
      RECT 70.176 67.691 71.864 67.759 ;
      RECT 70.222 67.645 71.91 67.713 ;
      RECT 70.268 67.599 71.956 67.667 ;
      RECT 70.314 67.553 72.002 67.621 ;
      RECT 70.36 67.507 72.048 67.575 ;
      RECT 70.406 67.461 72.094 67.529 ;
      RECT 70.452 67.415 72.14 67.483 ;
      RECT 70.498 67.369 72.186 67.437 ;
      RECT 70.544 67.323 72.232 67.391 ;
      RECT 70.59 67.277 72.278 67.345 ;
      RECT 70.636 67.231 72.324 67.299 ;
      RECT 70.682 67.185 72.37 67.253 ;
      RECT 70.728 67.139 72.416 67.207 ;
      RECT 70.774 67.093 72.462 67.161 ;
      RECT 70.82 67.047 72.508 67.115 ;
      RECT 70.866 67.001 72.554 67.069 ;
      RECT 70.912 66.955 72.6 67.023 ;
      RECT 70.958 66.909 72.646 66.977 ;
      RECT 71.004 66.863 72.692 66.931 ;
      RECT 71.05 66.817 72.738 66.885 ;
      RECT 71.096 66.771 72.784 66.839 ;
      RECT 71.142 66.725 72.83 66.793 ;
      RECT 71.188 66.679 72.876 66.747 ;
      RECT 71.234 66.633 72.922 66.701 ;
      RECT 71.28 66.587 72.968 66.655 ;
      RECT 71.326 66.541 73.014 66.609 ;
      RECT 71.372 66.495 73.06 66.563 ;
      RECT 71.418 66.449 73.106 66.517 ;
      RECT 71.464 66.403 73.152 66.471 ;
      RECT 71.51 66.357 73.198 66.425 ;
      RECT 71.556 66.311 73.244 66.379 ;
      RECT 71.602 66.265 73.29 66.333 ;
      RECT 71.648 66.219 73.336 66.287 ;
      RECT 71.694 66.173 73.382 66.241 ;
      RECT 71.74 66.127 73.428 66.195 ;
      RECT 71.786 66.081 73.474 66.149 ;
      RECT 71.832 66.035 73.52 66.103 ;
      RECT 71.878 65.989 73.566 66.057 ;
      RECT 71.924 65.943 73.612 66.011 ;
      RECT 71.97 65.897 73.658 65.965 ;
      RECT 72.016 65.851 73.704 65.919 ;
      RECT 72.062 65.805 73.75 65.873 ;
      RECT 72.108 65.759 73.796 65.827 ;
      RECT 72.154 65.713 73.842 65.781 ;
      RECT 72.2 65.667 73.888 65.735 ;
      RECT 72.246 65.621 73.934 65.689 ;
      RECT 72.292 65.575 73.98 65.643 ;
      RECT 72.338 65.529 74.026 65.597 ;
      RECT 72.384 65.483 74.072 65.551 ;
      RECT 72.43 65.437 74.118 65.505 ;
      RECT 72.476 65.391 74.164 65.459 ;
      RECT 72.522 65.345 74.21 65.413 ;
      RECT 72.568 65.299 74.256 65.367 ;
      RECT 72.614 65.253 74.302 65.321 ;
      RECT 72.66 65.207 74.348 65.275 ;
      RECT 72.706 65.161 74.394 65.229 ;
      RECT 72.752 65.115 74.44 65.183 ;
      RECT 72.798 65.069 74.486 65.137 ;
      RECT 72.844 65.023 74.532 65.091 ;
      RECT 72.89 64.977 74.578 65.045 ;
      RECT 72.936 64.931 74.624 64.999 ;
      RECT 72.982 64.885 74.67 64.953 ;
      RECT 73.028 64.839 74.716 64.907 ;
      RECT 73.074 64.793 74.762 64.861 ;
      RECT 73.12 64.747 74.808 64.815 ;
      RECT 73.166 64.701 74.854 64.769 ;
      RECT 73.212 64.655 74.9 64.723 ;
      RECT 73.258 64.609 74.946 64.677 ;
      RECT 73.304 64.563 74.992 64.631 ;
      RECT 73.35 64.517 75.038 64.585 ;
      RECT 73.396 64.471 75.084 64.539 ;
      RECT 73.442 64.425 75.13 64.493 ;
      RECT 73.488 64.379 75.176 64.447 ;
      RECT 73.534 64.333 75.222 64.401 ;
      RECT 73.58 64.287 75.268 64.355 ;
      RECT 73.626 64.241 75.314 64.309 ;
      RECT 73.672 64.195 75.36 64.263 ;
      RECT 73.718 64.149 75.406 64.217 ;
      RECT 73.764 64.103 75.452 64.171 ;
      RECT 73.81 64.057 75.498 64.125 ;
      RECT 73.856 64.011 75.544 64.079 ;
      RECT 73.902 63.965 75.59 64.033 ;
      RECT 73.948 63.919 75.636 63.987 ;
      RECT 73.994 63.873 75.682 63.941 ;
      RECT 74.04 63.827 75.728 63.895 ;
      RECT 74.086 63.781 75.774 63.849 ;
      RECT 74.132 63.735 75.82 63.803 ;
      RECT 74.178 63.689 75.866 63.757 ;
      RECT 74.224 63.643 75.912 63.711 ;
      RECT 74.27 63.597 75.958 63.665 ;
      RECT 74.316 63.551 76.004 63.619 ;
      RECT 74.362 63.505 76.05 63.573 ;
      RECT 74.408 63.459 76.096 63.527 ;
      RECT 74.454 63.413 76.142 63.481 ;
      RECT 74.5 63.367 76.188 63.435 ;
      RECT 74.546 63.321 76.234 63.389 ;
      RECT 74.592 63.275 76.28 63.343 ;
      RECT 74.638 63.229 76.326 63.297 ;
      RECT 74.684 63.183 76.372 63.251 ;
      RECT 74.73 63.137 76.418 63.205 ;
      RECT 74.776 63.091 76.464 63.159 ;
      RECT 74.822 63.045 76.51 63.113 ;
      RECT 74.868 62.999 76.556 63.067 ;
      RECT 74.914 62.953 76.602 63.021 ;
      RECT 76.57 61.308 76.602 63.021 ;
      RECT 74.96 62.907 76.648 62.975 ;
      RECT 76.595 61.272 76.648 62.975 ;
      RECT 75.006 62.861 76.694 62.929 ;
      RECT 76.641 61.226 76.694 62.929 ;
      RECT 75.052 62.815 76.74 62.883 ;
      RECT 76.687 61.18 76.74 62.883 ;
      RECT 75.098 62.769 76.786 62.837 ;
      RECT 76.733 61.134 76.786 62.837 ;
      RECT 75.144 62.723 76.832 62.791 ;
      RECT 76.779 61.088 76.832 62.791 ;
      RECT 75.19 62.677 76.878 62.745 ;
      RECT 76.825 61.042 76.878 62.745 ;
      RECT 75.236 62.631 76.924 62.699 ;
      RECT 76.871 60.996 76.924 62.699 ;
      RECT 75.282 62.585 76.97 62.653 ;
      RECT 76.917 60.95 76.97 62.653 ;
      RECT 75.328 62.539 77.016 62.607 ;
      RECT 76.963 60.904 77.016 62.607 ;
      RECT 75.374 62.493 77.062 62.561 ;
      RECT 77.009 60.858 77.062 62.561 ;
      RECT 75.42 62.447 77.108 62.515 ;
      RECT 77.055 60.812 77.108 62.515 ;
      RECT 75.466 62.401 77.154 62.469 ;
      RECT 77.101 60.766 77.154 62.469 ;
      RECT 75.512 62.355 77.2 62.423 ;
      RECT 77.147 60.72 77.2 62.423 ;
      RECT 75.558 62.309 77.246 62.377 ;
      RECT 77.193 60.674 77.246 62.377 ;
      RECT 75.604 62.263 77.292 62.331 ;
      RECT 77.239 60.628 77.292 62.331 ;
      RECT 75.65 62.217 77.338 62.285 ;
      RECT 77.285 60.582 77.338 62.285 ;
      RECT 75.696 62.171 77.384 62.239 ;
      RECT 77.331 60.536 77.384 62.239 ;
      RECT 75.742 62.125 77.43 62.193 ;
      RECT 77.377 60.49 77.43 62.193 ;
      RECT 75.788 62.079 77.476 62.147 ;
      RECT 77.423 60.444 77.476 62.147 ;
      RECT 75.834 62.033 77.522 62.101 ;
      RECT 77.469 60.398 77.522 62.101 ;
      RECT 75.88 61.987 77.568 62.055 ;
      RECT 77.515 60.352 77.568 62.055 ;
      RECT 75.926 61.941 77.614 62.009 ;
      RECT 77.561 60.306 77.614 62.009 ;
      RECT 75.972 61.895 77.66 61.963 ;
      RECT 77.607 60.26 77.66 61.963 ;
      RECT 76.018 61.849 77.706 61.917 ;
      RECT 77.653 60.214 77.706 61.917 ;
      RECT 76.064 61.803 77.752 61.871 ;
      RECT 77.699 60.168 77.752 61.871 ;
      RECT 76.11 61.757 77.798 61.825 ;
      RECT 77.745 60.122 77.798 61.825 ;
      RECT 76.156 61.711 77.844 61.779 ;
      RECT 77.791 60.076 77.844 61.779 ;
      RECT 76.202 61.665 77.89 61.733 ;
      RECT 77.837 60.03 77.89 61.733 ;
      RECT 76.248 61.619 77.936 61.687 ;
      RECT 77.883 59.984 77.936 61.687 ;
      RECT 76.294 61.573 77.982 61.641 ;
      RECT 77.929 59.938 77.982 61.641 ;
      RECT 76.34 61.527 78.028 61.595 ;
      RECT 77.975 59.892 78.028 61.595 ;
      RECT 76.386 61.481 78.074 61.549 ;
      RECT 78.021 59.846 78.074 61.549 ;
      RECT 76.432 61.435 78.12 61.503 ;
      RECT 78.067 59.8 78.12 61.503 ;
      RECT 76.478 61.389 78.166 61.457 ;
      RECT 78.113 59.754 78.166 61.457 ;
      RECT 76.524 61.343 78.212 61.411 ;
      RECT 78.159 59.708 78.212 61.411 ;
      RECT 78.205 59.662 78.258 61.365 ;
      RECT 78.251 59.616 78.304 61.319 ;
      RECT 78.297 59.57 78.35 61.273 ;
      RECT 78.343 59.524 78.396 61.227 ;
      RECT 78.389 59.478 78.442 61.181 ;
      RECT 78.435 59.432 78.488 61.135 ;
      RECT 78.481 59.386 78.534 61.089 ;
      RECT 78.527 59.34 78.58 61.043 ;
      RECT 78.573 59.294 78.626 60.997 ;
      RECT 78.619 59.248 78.672 60.951 ;
      RECT 78.665 59.202 78.718 60.905 ;
      RECT 78.711 59.156 78.764 60.859 ;
      RECT 78.757 59.11 78.81 60.813 ;
      RECT 78.803 59.064 78.856 60.767 ;
      RECT 78.849 59.018 78.902 60.721 ;
      RECT 78.895 58.972 78.948 60.675 ;
      RECT 78.941 58.926 78.994 60.629 ;
      RECT 78.987 58.88 79.04 60.583 ;
      RECT 79.033 58.834 79.086 60.537 ;
      RECT 79.079 58.788 79.132 60.491 ;
      RECT 79.125 58.742 79.178 60.445 ;
      RECT 79.171 58.696 79.224 60.399 ;
      RECT 79.217 58.65 79.27 60.353 ;
      RECT 79.263 58.604 79.316 60.307 ;
      RECT 79.309 58.558 79.362 60.261 ;
      RECT 79.355 58.512 79.408 60.215 ;
      RECT 79.401 58.466 79.454 60.169 ;
      RECT 79.447 58.42 79.5 60.123 ;
      RECT 79.493 58.374 79.546 60.077 ;
      RECT 79.539 58.328 79.592 60.031 ;
      RECT 79.585 58.282 79.638 59.985 ;
      RECT 79.631 58.236 79.684 59.939 ;
      RECT 79.677 58.19 79.73 59.893 ;
      RECT 79.723 58.144 79.776 59.847 ;
      RECT 79.769 58.098 79.822 59.801 ;
      RECT 79.815 58.052 79.868 59.755 ;
      RECT 79.861 58.006 79.914 59.709 ;
      RECT 79.907 57.96 79.96 59.663 ;
      RECT 79.953 57.914 80.006 59.617 ;
      RECT 79.999 57.868 80.052 59.571 ;
      RECT 80.045 57.822 80.098 59.525 ;
      RECT 80.091 57.776 80.144 59.479 ;
      RECT 80.137 57.73 80.19 59.433 ;
      RECT 80.183 57.684 80.236 59.387 ;
      RECT 80.229 57.638 80.282 59.341 ;
      RECT 80.275 57.592 80.328 59.295 ;
      RECT 80.321 57.546 80.374 59.249 ;
      RECT 80.367 57.5 80.42 59.203 ;
      RECT 80.413 57.454 80.466 59.157 ;
      RECT 80.459 57.408 80.512 59.111 ;
      RECT 80.505 57.362 80.558 59.065 ;
      RECT 80.551 57.316 80.604 59.019 ;
      RECT 80.597 57.27 80.65 58.973 ;
      RECT 80.643 57.224 80.696 58.927 ;
      RECT 80.689 57.178 80.742 58.881 ;
      RECT 80.735 57.132 80.788 58.835 ;
      RECT 80.781 57.086 80.834 58.789 ;
      RECT 80.827 57.04 80.88 58.743 ;
      RECT 80.873 56.994 80.926 58.697 ;
      RECT 80.919 56.948 80.972 58.651 ;
      RECT 80.965 56.902 81.018 58.605 ;
      RECT 81.011 56.856 81.064 58.559 ;
      RECT 81.057 56.81 81.11 58.513 ;
      RECT 81.103 56.764 81.156 58.467 ;
      RECT 81.149 56.718 81.202 58.421 ;
      RECT 81.195 56.672 81.248 58.375 ;
      RECT 81.241 56.626 81.294 58.329 ;
      RECT 81.287 56.58 81.34 58.283 ;
      RECT 81.333 56.534 81.386 58.237 ;
      RECT 81.379 56.488 81.432 58.191 ;
      RECT 81.425 56.442 81.478 58.145 ;
      RECT 81.471 56.396 81.524 58.099 ;
      RECT 81.517 56.352 81.57 58.053 ;
      RECT 81.56 56.33 81.616 58.007 ;
      RECT 81.56 56.33 81.662 57.961 ;
      RECT 81.56 56.33 81.708 57.915 ;
      RECT 81.56 56.33 81.754 57.869 ;
      RECT 81.56 56.33 81.8 57.823 ;
      RECT 81.56 56.33 81.846 57.777 ;
      RECT 81.56 56.33 81.892 57.731 ;
      RECT 81.56 56.33 81.938 57.685 ;
      RECT 81.56 56.33 81.984 57.639 ;
      RECT 81.56 56.33 82.03 57.593 ;
      RECT 81.56 56.33 82.076 57.547 ;
      RECT 81.56 56.33 82.122 57.501 ;
      RECT 81.56 56.33 82.168 57.455 ;
      RECT 81.56 56.33 82.214 57.409 ;
      RECT 81.56 56.33 82.26 57.363 ;
      RECT 81.56 56.33 82.306 57.317 ;
      RECT 81.56 56.33 82.352 57.271 ;
      RECT 81.56 56.33 82.398 57.225 ;
      RECT 81.56 56.33 82.43 57.186 ;
      RECT 81.56 56.33 110 57.17 ;
      RECT 63.83 85.547 68.17 110 ;
      RECT 63.83 85.547 68.216 88.012 ;
      RECT 63.83 85.547 68.262 87.966 ;
      RECT 63.83 85.547 68.308 87.92 ;
      RECT 63.83 85.547 68.354 87.874 ;
      RECT 63.83 85.547 68.4 87.828 ;
      RECT 63.83 85.547 68.446 87.782 ;
      RECT 63.83 85.547 68.492 87.736 ;
      RECT 63.83 85.547 68.538 87.69 ;
      RECT 63.83 85.547 68.584 87.644 ;
      RECT 63.83 85.547 68.63 87.598 ;
      RECT 63.83 85.547 68.676 87.552 ;
      RECT 63.83 85.547 68.722 87.506 ;
      RECT 63.83 85.547 68.768 87.46 ;
      RECT 63.83 85.547 68.814 87.414 ;
      RECT 63.83 85.547 68.86 87.368 ;
      RECT 63.83 85.547 68.906 87.322 ;
      RECT 63.83 85.547 68.952 87.276 ;
      RECT 63.83 85.547 68.998 87.23 ;
      RECT 63.83 85.547 69.044 87.184 ;
      RECT 63.83 85.547 69.09 87.138 ;
      RECT 63.83 85.547 69.136 87.092 ;
      RECT 63.83 85.547 69.182 87.046 ;
      RECT 63.83 85.547 69.228 87 ;
      RECT 63.83 85.547 69.274 86.954 ;
      RECT 63.83 85.547 69.32 86.908 ;
      RECT 63.83 85.547 69.366 86.862 ;
      RECT 63.83 85.547 69.412 86.816 ;
      RECT 63.83 85.547 69.458 86.77 ;
      RECT 63.83 85.547 69.504 86.724 ;
      RECT 63.83 85.547 69.55 86.678 ;
      RECT 63.83 85.547 69.596 86.632 ;
      RECT 63.83 85.547 69.642 86.586 ;
      RECT 63.83 85.547 69.688 86.54 ;
      RECT 63.83 85.547 69.734 86.494 ;
      RECT 63.83 85.547 69.78 86.448 ;
      RECT 63.83 85.547 69.826 86.402 ;
      RECT 63.83 85.547 69.872 86.356 ;
      RECT 63.83 85.547 69.918 86.31 ;
      RECT 63.83 85.547 69.964 86.264 ;
      RECT 63.83 85.547 70.01 86.218 ;
      RECT 63.83 85.547 70.056 86.172 ;
      RECT 63.83 85.547 70.102 86.126 ;
      RECT 63.83 85.547 70.148 86.08 ;
      RECT 63.83 85.547 70.194 86.034 ;
      RECT 63.83 85.547 70.24 85.988 ;
      RECT 63.83 85.547 70.286 85.942 ;
      RECT 63.83 85.547 70.332 85.896 ;
      RECT 63.83 85.547 70.378 85.85 ;
      RECT 63.83 85.547 70.424 85.804 ;
      RECT 63.83 85.547 70.47 85.758 ;
      RECT 63.83 85.547 70.516 85.712 ;
      RECT 63.83 85.547 70.562 85.666 ;
      RECT 63.83 85.547 70.608 85.62 ;
      RECT 63.876 85.501 70.654 85.574 ;
      RECT 70.592 78.785 70.654 85.574 ;
      RECT 63.922 85.455 70.7 85.528 ;
      RECT 70.638 78.739 70.7 85.528 ;
      RECT 63.968 85.409 70.746 85.482 ;
      RECT 70.684 78.693 70.746 85.482 ;
      RECT 64.014 85.363 70.792 85.436 ;
      RECT 70.73 78.647 70.792 85.436 ;
      RECT 64.06 85.317 70.838 85.39 ;
      RECT 70.776 78.601 70.838 85.39 ;
      RECT 64.106 85.271 70.884 85.344 ;
      RECT 70.822 78.555 70.884 85.344 ;
      RECT 64.152 85.225 70.93 85.298 ;
      RECT 70.868 78.509 70.93 85.298 ;
      RECT 64.198 85.179 70.976 85.252 ;
      RECT 70.914 78.463 70.976 85.252 ;
      RECT 64.244 85.133 71.022 85.206 ;
      RECT 70.96 78.417 71.022 85.206 ;
      RECT 64.29 85.087 71.068 85.16 ;
      RECT 71.006 78.371 71.068 85.16 ;
      RECT 64.336 85.041 71.114 85.114 ;
      RECT 71.052 78.325 71.114 85.114 ;
      RECT 64.382 84.995 71.16 85.068 ;
      RECT 71.098 78.279 71.16 85.068 ;
      RECT 64.428 84.949 71.206 85.022 ;
      RECT 71.144 78.233 71.206 85.022 ;
      RECT 64.474 84.903 71.252 84.976 ;
      RECT 71.19 78.187 71.252 84.976 ;
      RECT 64.52 84.857 71.298 84.93 ;
      RECT 71.236 78.141 71.298 84.93 ;
      RECT 64.566 84.811 71.344 84.884 ;
      RECT 71.282 78.095 71.344 84.884 ;
      RECT 64.612 84.765 71.39 84.838 ;
      RECT 71.328 78.049 71.39 84.838 ;
      RECT 64.658 84.719 71.436 84.792 ;
      RECT 71.374 78.003 71.436 84.792 ;
      RECT 64.704 84.673 71.482 84.746 ;
      RECT 71.42 77.957 71.482 84.746 ;
      RECT 64.75 84.627 71.528 84.7 ;
      RECT 71.466 77.911 71.528 84.7 ;
      RECT 64.796 84.581 71.574 84.654 ;
      RECT 71.512 77.865 71.574 84.654 ;
      RECT 64.842 84.535 71.62 84.608 ;
      RECT 71.558 77.819 71.62 84.608 ;
      RECT 64.888 84.489 71.666 84.562 ;
      RECT 71.604 77.773 71.666 84.562 ;
      RECT 64.934 84.443 71.712 84.516 ;
      RECT 71.65 77.727 71.712 84.516 ;
      RECT 64.98 84.397 71.758 84.47 ;
      RECT 71.696 77.681 71.758 84.47 ;
      RECT 65.026 84.351 71.804 84.424 ;
      RECT 71.742 77.635 71.804 84.424 ;
      RECT 65.072 84.305 71.85 84.378 ;
      RECT 71.788 77.589 71.85 84.378 ;
      RECT 65.118 84.259 71.896 84.332 ;
      RECT 71.834 77.543 71.896 84.332 ;
      RECT 65.164 84.213 71.942 84.286 ;
      RECT 71.88 77.497 71.942 84.286 ;
      RECT 65.21 84.167 71.988 84.24 ;
      RECT 71.926 77.451 71.988 84.24 ;
      RECT 65.256 84.121 72.034 84.194 ;
      RECT 71.972 77.405 72.034 84.194 ;
      RECT 65.302 84.075 72.08 84.148 ;
      RECT 72.018 77.359 72.08 84.148 ;
      RECT 65.348 84.029 72.126 84.102 ;
      RECT 72.064 77.313 72.126 84.102 ;
      RECT 65.394 83.983 72.172 84.056 ;
      RECT 72.11 77.267 72.172 84.056 ;
      RECT 65.44 83.937 72.218 84.01 ;
      RECT 72.156 77.221 72.218 84.01 ;
      RECT 65.486 83.891 72.264 83.964 ;
      RECT 72.202 77.175 72.264 83.964 ;
      RECT 65.532 83.845 72.31 83.918 ;
      RECT 72.248 77.129 72.31 83.918 ;
      RECT 65.578 83.799 72.356 83.872 ;
      RECT 72.294 77.083 72.356 83.872 ;
      RECT 65.624 83.753 72.402 83.826 ;
      RECT 72.34 77.037 72.402 83.826 ;
      RECT 65.67 83.707 72.448 83.78 ;
      RECT 72.386 76.991 72.448 83.78 ;
      RECT 65.716 83.661 72.494 83.734 ;
      RECT 72.432 76.945 72.494 83.734 ;
      RECT 65.762 83.615 72.54 83.688 ;
      RECT 72.478 76.899 72.54 83.688 ;
      RECT 65.808 83.569 72.586 83.642 ;
      RECT 72.524 76.853 72.586 83.642 ;
      RECT 65.854 83.523 72.632 83.596 ;
      RECT 72.57 76.807 72.632 83.596 ;
      RECT 65.9 83.477 72.678 83.55 ;
      RECT 72.616 76.761 72.678 83.55 ;
      RECT 65.946 83.431 72.724 83.504 ;
      RECT 72.662 76.715 72.724 83.504 ;
      RECT 65.992 83.385 72.77 83.458 ;
      RECT 72.708 76.669 72.77 83.458 ;
      RECT 66.038 83.339 72.816 83.412 ;
      RECT 72.754 76.623 72.816 83.412 ;
      RECT 66.084 83.293 72.862 83.366 ;
      RECT 72.8 76.577 72.862 83.366 ;
      RECT 66.13 83.247 72.908 83.32 ;
      RECT 72.846 76.531 72.908 83.32 ;
      RECT 66.176 83.201 72.954 83.274 ;
      RECT 72.892 76.485 72.954 83.274 ;
      RECT 66.222 83.155 73 83.228 ;
      RECT 72.938 76.439 73 83.228 ;
      RECT 66.268 83.109 73.046 83.182 ;
      RECT 72.984 76.393 73.046 83.182 ;
      RECT 66.314 83.063 73.092 83.136 ;
      RECT 73.03 76.347 73.092 83.136 ;
      RECT 66.36 83.017 73.138 83.09 ;
      RECT 73.076 76.301 73.138 83.09 ;
      RECT 66.406 82.971 73.184 83.044 ;
      RECT 73.122 76.255 73.184 83.044 ;
      RECT 66.452 82.925 73.23 82.998 ;
      RECT 73.168 76.209 73.23 82.998 ;
      RECT 66.498 82.879 73.276 82.952 ;
      RECT 73.214 76.163 73.276 82.952 ;
      RECT 66.544 82.833 73.322 82.906 ;
      RECT 73.26 76.117 73.322 82.906 ;
      RECT 66.59 82.787 73.368 82.86 ;
      RECT 73.306 76.071 73.368 82.86 ;
      RECT 66.636 82.741 73.414 82.814 ;
      RECT 73.352 76.025 73.414 82.814 ;
      RECT 66.682 82.695 73.46 82.768 ;
      RECT 73.398 75.979 73.46 82.768 ;
      RECT 66.728 82.649 73.506 82.722 ;
      RECT 73.444 75.933 73.506 82.722 ;
      RECT 66.774 82.603 73.552 82.676 ;
      RECT 73.49 75.887 73.552 82.676 ;
      RECT 66.82 82.557 73.598 82.63 ;
      RECT 73.536 75.841 73.598 82.63 ;
      RECT 66.866 82.511 73.644 82.584 ;
      RECT 73.582 75.795 73.644 82.584 ;
      RECT 66.912 82.465 73.69 82.538 ;
      RECT 73.628 75.749 73.69 82.538 ;
      RECT 66.958 82.419 73.736 82.492 ;
      RECT 73.674 75.703 73.736 82.492 ;
      RECT 67.004 82.373 73.782 82.446 ;
      RECT 73.72 75.657 73.782 82.446 ;
      RECT 67.05 82.327 73.828 82.4 ;
      RECT 73.766 75.611 73.828 82.4 ;
      RECT 67.096 82.281 73.874 82.354 ;
      RECT 73.812 75.565 73.874 82.354 ;
      RECT 67.142 82.235 73.92 82.308 ;
      RECT 73.858 75.519 73.92 82.308 ;
      RECT 67.188 82.189 73.966 82.262 ;
      RECT 73.904 75.473 73.966 82.262 ;
      RECT 67.234 82.143 74.012 82.216 ;
      RECT 73.95 75.427 74.012 82.216 ;
      RECT 67.28 82.097 74.058 82.17 ;
      RECT 73.996 75.381 74.058 82.17 ;
      RECT 67.326 82.051 74.104 82.124 ;
      RECT 74.042 75.335 74.104 82.124 ;
      RECT 67.372 82.005 74.15 82.078 ;
      RECT 74.088 75.289 74.15 82.078 ;
      RECT 67.418 81.959 74.196 82.032 ;
      RECT 74.134 75.243 74.196 82.032 ;
      RECT 67.464 81.913 74.242 81.986 ;
      RECT 74.18 75.197 74.242 81.986 ;
      RECT 67.51 81.867 74.288 81.94 ;
      RECT 74.226 75.151 74.288 81.94 ;
      RECT 67.556 81.821 74.334 81.894 ;
      RECT 74.272 75.105 74.334 81.894 ;
      RECT 67.602 81.775 74.38 81.848 ;
      RECT 74.318 75.059 74.38 81.848 ;
      RECT 67.648 81.729 74.426 81.802 ;
      RECT 74.364 75.013 74.426 81.802 ;
      RECT 67.694 81.683 74.472 81.756 ;
      RECT 74.41 74.967 74.472 81.756 ;
      RECT 67.74 81.637 74.518 81.71 ;
      RECT 74.456 74.921 74.518 81.71 ;
      RECT 67.786 81.591 74.564 81.664 ;
      RECT 74.502 74.875 74.564 81.664 ;
      RECT 67.832 81.545 74.61 81.618 ;
      RECT 74.548 74.829 74.61 81.618 ;
      RECT 67.878 81.499 74.656 81.572 ;
      RECT 74.594 74.783 74.656 81.572 ;
      RECT 67.924 81.453 74.702 81.526 ;
      RECT 74.64 74.737 74.702 81.526 ;
      RECT 67.97 81.407 74.748 81.48 ;
      RECT 74.686 74.691 74.748 81.48 ;
      RECT 68.016 81.361 74.794 81.434 ;
      RECT 74.732 74.645 74.794 81.434 ;
      RECT 68.062 81.315 74.84 81.388 ;
      RECT 74.778 74.599 74.84 81.388 ;
      RECT 68.108 81.269 74.886 81.342 ;
      RECT 74.824 74.553 74.886 81.342 ;
      RECT 68.154 81.223 74.932 81.296 ;
      RECT 74.87 74.507 74.932 81.296 ;
      RECT 68.2 81.177 74.978 81.25 ;
      RECT 74.916 74.461 74.978 81.25 ;
      RECT 68.246 81.131 75.024 81.204 ;
      RECT 74.962 74.415 75.024 81.204 ;
      RECT 68.292 81.085 75.07 81.158 ;
      RECT 75.008 74.369 75.07 81.158 ;
      RECT 68.338 81.039 75.116 81.112 ;
      RECT 75.054 74.323 75.116 81.112 ;
      RECT 68.384 80.993 75.162 81.066 ;
      RECT 75.1 74.277 75.162 81.066 ;
      RECT 68.43 80.947 75.208 81.02 ;
      RECT 75.146 74.231 75.208 81.02 ;
      RECT 68.476 80.901 75.254 80.974 ;
      RECT 75.192 74.185 75.254 80.974 ;
      RECT 68.522 80.855 75.3 80.928 ;
      RECT 75.238 74.139 75.3 80.928 ;
      RECT 68.568 80.809 75.346 80.882 ;
      RECT 75.284 74.093 75.346 80.882 ;
      RECT 68.614 80.763 75.392 80.836 ;
      RECT 75.33 74.047 75.392 80.836 ;
      RECT 68.66 80.717 75.438 80.79 ;
      RECT 75.376 74.001 75.438 80.79 ;
      RECT 68.706 80.671 75.484 80.744 ;
      RECT 75.422 73.955 75.484 80.744 ;
      RECT 68.752 80.625 75.53 80.698 ;
      RECT 75.468 73.909 75.53 80.698 ;
      RECT 68.798 80.579 75.576 80.652 ;
      RECT 75.514 73.863 75.576 80.652 ;
      RECT 68.844 80.533 75.622 80.606 ;
      RECT 75.56 73.817 75.622 80.606 ;
      RECT 68.89 80.487 75.668 80.56 ;
      RECT 75.606 73.771 75.668 80.56 ;
      RECT 68.936 80.441 75.714 80.514 ;
      RECT 75.652 73.725 75.714 80.514 ;
      RECT 68.982 80.395 75.76 80.468 ;
      RECT 75.698 73.679 75.76 80.468 ;
      RECT 69.028 80.349 75.806 80.422 ;
      RECT 75.744 73.633 75.806 80.422 ;
      RECT 69.074 80.303 75.852 80.376 ;
      RECT 75.79 73.587 75.852 80.376 ;
      RECT 69.12 80.257 75.898 80.33 ;
      RECT 75.836 73.541 75.898 80.33 ;
      RECT 69.166 80.211 75.944 80.284 ;
      RECT 75.882 73.495 75.944 80.284 ;
      RECT 69.212 80.165 75.99 80.238 ;
      RECT 75.928 73.449 75.99 80.238 ;
      RECT 69.258 80.119 76.036 80.192 ;
      RECT 75.974 73.403 76.036 80.192 ;
      RECT 69.304 80.073 76.082 80.146 ;
      RECT 76.02 73.357 76.082 80.146 ;
      RECT 69.35 80.027 76.128 80.1 ;
      RECT 76.066 73.311 76.128 80.1 ;
      RECT 69.396 79.981 76.174 80.054 ;
      RECT 76.112 73.265 76.174 80.054 ;
      RECT 69.442 79.935 76.22 80.008 ;
      RECT 76.158 73.219 76.22 80.008 ;
      RECT 69.488 79.889 76.266 79.962 ;
      RECT 76.204 73.173 76.266 79.962 ;
      RECT 69.534 79.843 76.312 79.916 ;
      RECT 76.25 73.127 76.312 79.916 ;
      RECT 69.58 79.797 76.358 79.87 ;
      RECT 76.296 73.081 76.358 79.87 ;
      RECT 69.626 79.751 76.404 79.824 ;
      RECT 76.342 73.035 76.404 79.824 ;
      RECT 69.672 79.705 76.45 79.778 ;
      RECT 76.388 72.989 76.45 79.778 ;
      RECT 69.718 79.659 76.496 79.732 ;
      RECT 76.434 72.943 76.496 79.732 ;
      RECT 69.764 79.613 76.542 79.686 ;
      RECT 76.48 72.897 76.542 79.686 ;
      RECT 69.81 79.567 76.588 79.64 ;
      RECT 76.526 72.851 76.588 79.64 ;
      RECT 69.856 79.521 76.634 79.594 ;
      RECT 76.572 72.805 76.634 79.594 ;
      RECT 69.902 79.475 76.67 79.553 ;
      RECT 76.618 72.759 76.67 79.553 ;
      RECT 69.948 79.429 76.716 79.512 ;
      RECT 76.664 72.713 76.716 79.512 ;
      RECT 69.994 79.383 76.762 79.466 ;
      RECT 76.71 72.667 76.762 79.466 ;
      RECT 70.04 79.337 76.808 79.42 ;
      RECT 76.756 72.621 76.808 79.42 ;
      RECT 70.086 79.291 76.854 79.374 ;
      RECT 76.802 72.575 76.854 79.374 ;
      RECT 70.132 79.245 76.9 79.328 ;
      RECT 76.848 72.529 76.9 79.328 ;
      RECT 70.178 79.199 76.946 79.282 ;
      RECT 76.894 72.483 76.946 79.282 ;
      RECT 70.224 79.153 76.992 79.236 ;
      RECT 76.94 72.437 76.992 79.236 ;
      RECT 70.27 79.107 77.038 79.19 ;
      RECT 76.986 72.391 77.038 79.19 ;
      RECT 70.316 79.061 77.084 79.144 ;
      RECT 77.032 72.345 77.084 79.144 ;
      RECT 70.362 79.015 77.13 79.098 ;
      RECT 77.078 72.299 77.13 79.098 ;
      RECT 70.408 78.969 77.176 79.052 ;
      RECT 77.124 72.253 77.176 79.052 ;
      RECT 70.454 78.923 77.222 79.006 ;
      RECT 77.17 72.207 77.222 79.006 ;
      RECT 70.5 78.877 77.268 78.96 ;
      RECT 77.216 72.161 77.268 78.96 ;
      RECT 70.546 78.831 77.314 78.914 ;
      RECT 77.262 72.115 77.314 78.914 ;
      RECT 77.308 72.069 77.36 78.868 ;
      RECT 77.354 72.023 77.406 78.822 ;
      RECT 77.4 71.977 77.452 78.776 ;
      RECT 77.446 71.931 77.498 78.73 ;
      RECT 77.492 71.885 77.544 78.684 ;
      RECT 77.538 71.839 77.59 78.638 ;
      RECT 77.584 71.793 77.636 78.592 ;
      RECT 77.63 71.747 77.682 78.546 ;
      RECT 77.676 71.701 77.728 78.5 ;
      RECT 77.722 71.655 77.774 78.454 ;
      RECT 77.768 71.609 77.82 78.408 ;
      RECT 77.814 71.563 77.866 78.362 ;
      RECT 77.86 71.517 77.912 78.316 ;
      RECT 77.906 71.471 77.958 78.27 ;
      RECT 77.952 71.425 78.004 78.224 ;
      RECT 77.998 71.379 78.05 78.178 ;
      RECT 78.044 71.333 78.096 78.132 ;
      RECT 78.09 71.287 78.142 78.086 ;
      RECT 78.136 71.241 78.188 78.04 ;
      RECT 78.182 71.195 78.234 77.994 ;
      RECT 78.228 71.149 78.28 77.948 ;
      RECT 78.274 71.103 78.326 77.902 ;
      RECT 78.32 71.057 78.372 77.856 ;
      RECT 78.366 71.011 78.418 77.81 ;
      RECT 78.412 70.965 78.464 77.764 ;
      RECT 78.458 70.919 78.51 77.718 ;
      RECT 78.504 70.873 78.556 77.672 ;
      RECT 78.55 70.827 78.602 77.626 ;
      RECT 78.596 70.781 78.648 77.58 ;
      RECT 78.642 70.735 78.694 77.534 ;
      RECT 78.688 70.689 78.74 77.488 ;
      RECT 78.734 70.643 78.786 77.442 ;
      RECT 78.78 70.597 78.832 77.396 ;
      RECT 78.826 70.551 78.878 77.35 ;
      RECT 78.872 70.505 78.924 77.304 ;
      RECT 78.918 70.459 78.97 77.258 ;
      RECT 78.964 70.413 79.016 77.212 ;
      RECT 79.01 70.367 79.062 77.166 ;
      RECT 79.056 70.321 79.108 77.12 ;
      RECT 79.102 70.275 79.154 77.074 ;
      RECT 79.148 70.229 79.2 77.028 ;
      RECT 79.194 70.183 79.246 76.982 ;
      RECT 79.24 70.137 79.292 76.936 ;
      RECT 79.286 70.091 79.338 76.89 ;
      RECT 79.332 70.045 79.384 76.844 ;
      RECT 79.378 69.999 79.43 76.798 ;
      RECT 79.424 69.953 79.476 76.752 ;
      RECT 79.47 69.907 79.522 76.706 ;
      RECT 79.516 69.861 79.568 76.66 ;
      RECT 79.562 69.815 79.614 76.614 ;
      RECT 79.608 69.769 79.66 76.568 ;
      RECT 79.654 69.723 79.706 76.522 ;
      RECT 79.7 69.677 79.752 76.476 ;
      RECT 79.746 69.631 79.798 76.43 ;
      RECT 79.792 69.585 79.844 76.384 ;
      RECT 79.838 69.539 79.89 76.338 ;
      RECT 79.884 69.493 79.936 76.292 ;
      RECT 79.93 69.447 79.982 76.246 ;
      RECT 79.976 69.401 80.028 76.2 ;
      RECT 80.022 69.355 80.074 76.154 ;
      RECT 80.068 69.309 80.12 76.108 ;
      RECT 80.114 69.263 80.166 76.062 ;
      RECT 80.16 69.217 80.212 76.016 ;
      RECT 80.206 69.171 80.258 75.97 ;
      RECT 80.252 69.125 80.304 75.924 ;
      RECT 80.298 69.079 80.35 75.878 ;
      RECT 80.344 69.033 80.396 75.832 ;
      RECT 80.39 68.987 80.442 75.786 ;
      RECT 80.436 68.941 80.488 75.74 ;
      RECT 80.482 68.895 80.534 75.694 ;
      RECT 80.528 68.849 80.58 75.648 ;
      RECT 80.574 68.803 80.626 75.602 ;
      RECT 80.62 68.757 80.672 75.556 ;
      RECT 80.666 68.711 80.718 75.51 ;
      RECT 80.712 68.665 80.764 75.464 ;
      RECT 80.758 68.619 80.81 75.418 ;
      RECT 80.804 68.573 80.856 75.372 ;
      RECT 80.85 68.527 80.902 75.326 ;
      RECT 80.896 68.481 80.948 75.28 ;
      RECT 80.942 68.435 80.994 75.234 ;
      RECT 80.988 68.389 81.04 75.188 ;
      RECT 81.034 68.343 81.086 75.142 ;
      RECT 81.08 68.297 81.132 75.096 ;
      RECT 81.126 68.251 81.178 75.05 ;
      RECT 81.172 68.205 81.224 75.004 ;
      RECT 81.218 68.159 81.27 74.958 ;
      RECT 81.264 68.113 81.316 74.912 ;
      RECT 81.31 68.067 81.362 74.866 ;
      RECT 81.356 68.021 81.408 74.82 ;
      RECT 81.402 67.975 81.454 74.774 ;
      RECT 81.448 67.929 81.5 74.728 ;
      RECT 81.494 67.883 81.546 74.682 ;
      RECT 81.54 67.837 81.592 74.636 ;
      RECT 81.586 67.791 81.638 74.59 ;
      RECT 81.632 67.745 81.684 74.544 ;
      RECT 81.678 67.699 81.73 74.498 ;
      RECT 81.724 67.653 81.776 74.452 ;
      RECT 81.77 67.607 81.822 74.406 ;
      RECT 81.816 67.561 81.868 74.36 ;
      RECT 81.862 67.515 81.914 74.314 ;
      RECT 81.908 67.469 81.96 74.268 ;
      RECT 81.954 67.423 82.006 74.222 ;
      RECT 82 67.377 82.052 74.176 ;
      RECT 82.046 67.331 82.098 74.13 ;
      RECT 82.092 67.285 82.144 74.084 ;
      RECT 82.138 67.239 82.19 74.038 ;
      RECT 82.184 67.193 82.236 73.992 ;
      RECT 82.23 67.147 82.282 73.946 ;
      RECT 82.276 67.101 82.328 73.9 ;
      RECT 82.322 67.055 82.374 73.854 ;
      RECT 82.368 67.009 82.42 73.808 ;
      RECT 82.414 66.963 82.466 73.762 ;
      RECT 82.46 66.917 82.512 73.716 ;
      RECT 82.506 66.871 82.558 73.67 ;
      RECT 82.552 66.825 82.604 73.624 ;
      RECT 82.598 66.779 82.65 73.578 ;
      RECT 82.644 66.733 82.696 73.532 ;
      RECT 82.69 66.687 82.742 73.486 ;
      RECT 82.736 66.641 82.788 73.44 ;
      RECT 82.782 66.595 82.834 73.394 ;
      RECT 82.828 66.549 82.88 73.348 ;
      RECT 82.874 66.503 82.926 73.302 ;
      RECT 82.92 66.457 82.972 73.256 ;
      RECT 82.966 66.411 83.018 73.21 ;
      RECT 83.012 66.365 83.064 73.164 ;
      RECT 83.058 66.326 83.11 73.118 ;
      RECT 83.09 66.287 83.156 73.072 ;
      RECT 83.136 66.241 83.202 73.026 ;
      RECT 83.182 66.195 83.248 72.98 ;
      RECT 83.228 66.149 83.294 72.934 ;
      RECT 83.274 66.103 83.34 72.888 ;
      RECT 83.32 66.057 83.386 72.842 ;
      RECT 83.366 66.011 83.432 72.796 ;
      RECT 83.412 65.965 83.478 72.75 ;
      RECT 83.458 65.919 83.524 72.704 ;
      RECT 83.504 65.873 83.57 72.658 ;
      RECT 83.55 65.827 83.616 72.612 ;
      RECT 83.596 65.781 83.662 72.566 ;
      RECT 83.642 65.735 83.708 72.52 ;
      RECT 83.688 65.689 83.754 72.474 ;
      RECT 83.734 65.643 83.8 72.428 ;
      RECT 83.78 65.597 83.846 72.382 ;
      RECT 83.826 65.551 83.892 72.336 ;
      RECT 83.872 65.505 83.938 72.29 ;
      RECT 83.918 65.459 83.984 72.244 ;
      RECT 83.964 65.413 84.03 72.198 ;
      RECT 84.01 65.367 84.076 72.152 ;
      RECT 84.056 65.321 84.122 72.106 ;
      RECT 84.102 65.275 84.168 72.06 ;
      RECT 84.148 65.229 84.214 72.014 ;
      RECT 84.194 65.183 84.26 71.968 ;
      RECT 84.24 65.137 84.306 71.922 ;
      RECT 84.286 65.091 84.352 71.876 ;
      RECT 84.332 65.045 84.398 71.83 ;
      RECT 84.378 64.999 84.444 71.784 ;
      RECT 84.424 64.953 84.49 71.738 ;
      RECT 84.47 64.907 84.536 71.692 ;
      RECT 84.516 64.861 84.582 71.646 ;
      RECT 84.562 64.815 84.628 71.6 ;
      RECT 84.608 64.769 84.674 71.554 ;
      RECT 84.654 64.723 84.72 71.508 ;
      RECT 84.7 64.677 84.766 71.462 ;
      RECT 84.746 64.631 84.812 71.416 ;
      RECT 84.792 64.585 84.858 71.37 ;
      RECT 84.838 64.539 84.904 71.324 ;
      RECT 84.884 64.493 84.95 71.278 ;
      RECT 84.93 64.447 84.996 71.232 ;
      RECT 84.976 64.401 85.042 71.186 ;
      RECT 85.022 64.355 85.088 71.14 ;
      RECT 85.068 64.309 85.134 71.094 ;
      RECT 85.114 64.263 85.18 71.048 ;
      RECT 85.16 64.217 85.226 71.002 ;
      RECT 85.206 64.171 85.272 70.956 ;
      RECT 85.252 64.125 85.318 70.91 ;
      RECT 85.298 64.079 85.364 70.864 ;
      RECT 85.344 64.033 85.41 70.818 ;
      RECT 85.39 63.987 85.456 70.772 ;
      RECT 85.436 63.941 85.502 70.726 ;
      RECT 85.482 63.895 85.548 70.68 ;
      RECT 85.528 63.851 85.594 70.634 ;
      RECT 85.57 63.83 85.64 70.588 ;
      RECT 85.57 63.83 85.686 70.542 ;
      RECT 85.57 63.83 85.732 70.496 ;
      RECT 85.57 63.83 85.778 70.45 ;
      RECT 85.57 63.83 85.824 70.404 ;
      RECT 85.57 63.83 85.87 70.358 ;
      RECT 85.57 63.83 85.916 70.312 ;
      RECT 85.57 63.83 85.962 70.266 ;
      RECT 85.57 63.83 86.008 70.22 ;
      RECT 85.57 63.83 86.054 70.174 ;
      RECT 85.57 63.83 86.1 70.128 ;
      RECT 85.57 63.83 86.146 70.082 ;
      RECT 85.57 63.83 86.192 70.036 ;
      RECT 85.57 63.83 86.238 69.99 ;
      RECT 85.57 63.83 86.284 69.944 ;
      RECT 85.57 63.83 86.33 69.898 ;
      RECT 85.57 63.83 86.376 69.852 ;
      RECT 85.57 63.83 86.422 69.806 ;
      RECT 85.57 63.83 86.468 69.76 ;
      RECT 85.57 63.83 86.514 69.714 ;
      RECT 85.57 63.83 86.56 69.668 ;
      RECT 85.57 63.83 86.606 69.622 ;
      RECT 85.57 63.83 86.652 69.576 ;
      RECT 85.57 63.83 86.698 69.53 ;
      RECT 85.57 63.83 86.744 69.484 ;
      RECT 85.57 63.83 86.79 69.438 ;
      RECT 85.57 63.83 86.836 69.392 ;
      RECT 85.57 63.83 86.882 69.346 ;
      RECT 85.57 63.83 86.928 69.3 ;
      RECT 85.57 63.83 86.974 69.254 ;
      RECT 85.57 63.83 87.02 69.208 ;
      RECT 85.57 63.83 87.066 69.162 ;
      RECT 85.57 63.83 87.112 69.116 ;
      RECT 85.57 63.83 87.158 69.07 ;
      RECT 85.57 63.83 87.204 69.024 ;
      RECT 85.57 63.83 87.25 68.978 ;
      RECT 85.57 63.83 87.296 68.932 ;
      RECT 85.57 63.83 87.342 68.886 ;
      RECT 85.57 63.83 87.388 68.84 ;
      RECT 85.57 63.83 87.434 68.794 ;
      RECT 85.57 63.83 87.48 68.748 ;
      RECT 85.57 63.83 87.526 68.702 ;
      RECT 85.57 63.83 87.572 68.656 ;
      RECT 85.57 63.83 87.618 68.61 ;
      RECT 85.57 63.83 87.664 68.564 ;
      RECT 85.57 63.83 87.71 68.518 ;
      RECT 85.57 63.83 87.756 68.472 ;
      RECT 85.57 63.83 87.802 68.426 ;
      RECT 85.57 63.83 87.848 68.38 ;
      RECT 85.57 63.83 87.894 68.334 ;
      RECT 85.57 63.83 87.94 68.288 ;
      RECT 85.57 63.83 87.986 68.242 ;
      RECT 81.218 68.159 88.032 68.196 ;
      RECT 81.218 68.159 88.035 68.171 ;
      RECT 85.57 63.83 110 68.17 ;
      RECT 77.33 92.192 78.17 110 ;
      RECT 77.376 92.146 78.17 110 ;
      RECT 77.422 92.1 78.17 110 ;
      RECT 77.468 92.054 78.216 92.117 ;
      RECT 77.514 92.008 78.262 92.071 ;
      RECT 77.56 91.962 78.308 92.025 ;
      RECT 77.606 91.916 78.354 91.979 ;
      RECT 77.652 91.87 78.4 91.933 ;
      RECT 77.698 91.824 78.446 91.887 ;
      RECT 77.744 91.778 78.492 91.841 ;
      RECT 77.79 91.732 78.538 91.795 ;
      RECT 77.836 91.686 78.584 91.749 ;
      RECT 77.882 91.64 78.63 91.703 ;
      RECT 77.928 91.594 78.676 91.657 ;
      RECT 77.974 91.548 78.722 91.611 ;
      RECT 78.02 91.502 78.768 91.565 ;
      RECT 78.066 91.456 78.814 91.519 ;
      RECT 78.112 91.41 78.86 91.473 ;
      RECT 78.158 91.364 78.906 91.427 ;
      RECT 78.204 91.318 78.952 91.381 ;
      RECT 78.25 91.272 78.998 91.335 ;
      RECT 78.296 91.226 79.044 91.289 ;
      RECT 78.342 91.18 79.09 91.243 ;
      RECT 78.388 91.134 79.136 91.197 ;
      RECT 78.434 91.088 79.182 91.151 ;
      RECT 78.48 91.042 79.228 91.105 ;
      RECT 78.526 90.996 79.274 91.059 ;
      RECT 78.572 90.95 79.32 91.013 ;
      RECT 78.618 90.904 79.366 90.967 ;
      RECT 78.664 90.858 79.412 90.921 ;
      RECT 78.71 90.812 79.458 90.875 ;
      RECT 78.756 90.766 79.504 90.829 ;
      RECT 78.802 90.72 79.55 90.783 ;
      RECT 78.848 90.674 79.596 90.737 ;
      RECT 78.894 90.628 79.642 90.691 ;
      RECT 78.94 90.582 79.688 90.645 ;
      RECT 78.986 90.536 79.734 90.599 ;
      RECT 79.032 90.49 79.78 90.553 ;
      RECT 79.078 90.444 79.826 90.507 ;
      RECT 79.124 90.398 79.872 90.461 ;
      RECT 79.17 90.352 79.918 90.415 ;
      RECT 79.216 90.306 79.964 90.369 ;
      RECT 79.262 90.26 80.01 90.323 ;
      RECT 79.308 90.214 80.056 90.277 ;
      RECT 79.354 90.168 80.102 90.231 ;
      RECT 79.4 90.122 80.148 90.185 ;
      RECT 79.446 90.076 80.194 90.139 ;
      RECT 79.492 90.03 80.24 90.093 ;
      RECT 79.538 89.984 80.286 90.047 ;
      RECT 79.584 89.938 80.332 90.001 ;
      RECT 79.63 89.892 80.378 89.955 ;
      RECT 79.676 89.846 80.424 89.909 ;
      RECT 79.722 89.8 80.47 89.863 ;
      RECT 79.768 89.754 80.516 89.817 ;
      RECT 79.814 89.708 80.562 89.771 ;
      RECT 79.86 89.662 80.608 89.725 ;
      RECT 79.906 89.616 80.654 89.679 ;
      RECT 79.952 89.57 80.7 89.633 ;
      RECT 79.998 89.524 80.746 89.587 ;
      RECT 80.044 89.478 80.792 89.541 ;
      RECT 80.09 89.432 80.838 89.495 ;
      RECT 80.136 89.386 80.884 89.449 ;
      RECT 80.182 89.34 80.93 89.403 ;
      RECT 80.228 89.294 80.976 89.357 ;
      RECT 80.274 89.248 81.022 89.311 ;
      RECT 80.32 89.202 81.068 89.265 ;
      RECT 80.366 89.156 81.114 89.219 ;
      RECT 80.412 89.11 81.16 89.173 ;
      RECT 80.458 89.064 81.206 89.127 ;
      RECT 80.504 89.018 81.252 89.081 ;
      RECT 80.55 88.972 81.298 89.035 ;
      RECT 80.596 88.926 81.344 88.989 ;
      RECT 80.642 88.88 81.39 88.943 ;
      RECT 80.688 88.834 81.436 88.897 ;
      RECT 80.734 88.788 81.482 88.851 ;
      RECT 80.78 88.742 81.528 88.805 ;
      RECT 80.826 88.696 81.574 88.759 ;
      RECT 80.872 88.65 81.62 88.713 ;
      RECT 80.918 88.604 81.666 88.667 ;
      RECT 80.964 88.558 81.712 88.621 ;
      RECT 81.01 88.512 81.758 88.575 ;
      RECT 81.056 88.466 81.804 88.529 ;
      RECT 81.102 88.42 81.85 88.483 ;
      RECT 81.148 88.374 81.896 88.437 ;
      RECT 81.194 88.328 81.942 88.391 ;
      RECT 81.24 88.282 81.988 88.345 ;
      RECT 81.286 88.236 82.034 88.299 ;
      RECT 81.332 88.19 82.08 88.253 ;
      RECT 81.378 88.144 82.126 88.207 ;
      RECT 81.424 88.098 82.172 88.161 ;
      RECT 81.47 88.052 82.218 88.115 ;
      RECT 81.516 88.006 82.264 88.069 ;
      RECT 81.562 87.96 82.31 88.023 ;
      RECT 81.608 87.914 82.356 87.977 ;
      RECT 81.654 87.868 82.402 87.931 ;
      RECT 81.7 87.822 82.448 87.885 ;
      RECT 81.746 87.776 82.494 87.839 ;
      RECT 81.792 87.73 82.54 87.793 ;
      RECT 81.838 87.684 82.586 87.747 ;
      RECT 81.884 87.638 82.632 87.701 ;
      RECT 81.93 87.592 82.678 87.655 ;
      RECT 81.976 87.546 82.724 87.609 ;
      RECT 82.022 87.5 82.77 87.563 ;
      RECT 82.068 87.454 82.816 87.517 ;
      RECT 82.114 87.408 82.862 87.471 ;
      RECT 82.16 87.362 82.908 87.425 ;
      RECT 82.206 87.316 82.954 87.379 ;
      RECT 82.252 87.27 83 87.333 ;
      RECT 82.298 87.224 83.046 87.287 ;
      RECT 82.344 87.178 83.092 87.241 ;
      RECT 82.39 87.132 83.138 87.195 ;
      RECT 82.436 87.086 83.184 87.149 ;
      RECT 82.482 87.04 83.23 87.103 ;
      RECT 82.528 86.994 83.276 87.057 ;
      RECT 82.574 86.948 83.322 87.011 ;
      RECT 82.62 86.902 83.368 86.965 ;
      RECT 82.666 86.856 83.414 86.919 ;
      RECT 82.712 86.81 83.46 86.873 ;
      RECT 82.758 86.764 83.506 86.827 ;
      RECT 82.804 86.718 83.552 86.781 ;
      RECT 82.85 86.672 83.598 86.735 ;
      RECT 82.896 86.626 83.644 86.689 ;
      RECT 82.942 86.58 83.69 86.643 ;
      RECT 82.988 86.534 83.736 86.597 ;
      RECT 83.034 86.488 83.782 86.551 ;
      RECT 83.08 86.442 83.828 86.505 ;
      RECT 83.126 86.396 83.874 86.459 ;
      RECT 83.172 86.35 83.92 86.413 ;
      RECT 83.218 86.304 83.966 86.367 ;
      RECT 83.264 86.258 84.012 86.321 ;
      RECT 83.31 86.212 84.058 86.275 ;
      RECT 83.356 86.166 84.104 86.229 ;
      RECT 83.402 86.12 84.15 86.183 ;
      RECT 83.448 86.074 84.196 86.137 ;
      RECT 83.494 86.028 84.242 86.091 ;
      RECT 83.54 85.982 84.288 86.045 ;
      RECT 83.586 85.936 84.334 85.999 ;
      RECT 83.632 85.89 84.38 85.953 ;
      RECT 83.678 85.844 84.426 85.907 ;
      RECT 83.724 85.798 84.472 85.861 ;
      RECT 83.77 85.752 84.518 85.815 ;
      RECT 83.816 85.706 84.564 85.769 ;
      RECT 83.862 85.66 84.61 85.723 ;
      RECT 83.908 85.614 84.656 85.677 ;
      RECT 83.954 85.568 84.702 85.631 ;
      RECT 84 85.522 84.748 85.585 ;
      RECT 84.046 85.476 84.794 85.539 ;
      RECT 84.092 85.43 84.84 85.493 ;
      RECT 84.138 85.384 84.886 85.447 ;
      RECT 84.184 85.338 84.932 85.401 ;
      RECT 84.23 85.292 84.978 85.355 ;
      RECT 84.276 85.246 85.024 85.309 ;
      RECT 84.322 85.2 85.07 85.263 ;
      RECT 84.368 85.154 85.116 85.217 ;
      RECT 84.414 85.108 85.162 85.171 ;
      RECT 84.46 85.062 85.208 85.125 ;
      RECT 84.506 85.016 85.254 85.079 ;
      RECT 84.552 84.97 85.3 85.033 ;
      RECT 84.598 84.924 85.346 84.987 ;
      RECT 84.644 84.878 85.392 84.941 ;
      RECT 84.69 84.832 85.438 84.895 ;
      RECT 84.736 84.786 85.484 84.849 ;
      RECT 84.782 84.74 85.53 84.803 ;
      RECT 84.828 84.694 85.576 84.757 ;
      RECT 84.874 84.648 85.622 84.711 ;
      RECT 84.92 84.602 85.668 84.665 ;
      RECT 84.966 84.556 85.714 84.619 ;
      RECT 85.012 84.51 85.76 84.573 ;
      RECT 85.058 84.464 85.806 84.527 ;
      RECT 85.104 84.418 85.852 84.481 ;
      RECT 85.15 84.372 85.898 84.435 ;
      RECT 85.196 84.326 85.944 84.389 ;
      RECT 85.242 84.28 85.99 84.343 ;
      RECT 85.288 84.234 86.036 84.297 ;
      RECT 85.334 84.188 86.082 84.251 ;
      RECT 85.38 84.142 86.128 84.205 ;
      RECT 85.426 84.096 86.174 84.159 ;
      RECT 85.472 84.05 86.22 84.113 ;
      RECT 85.518 84.004 86.266 84.067 ;
      RECT 85.564 83.958 86.312 84.021 ;
      RECT 85.61 83.912 86.358 83.975 ;
      RECT 85.656 83.866 86.404 83.929 ;
      RECT 85.702 83.82 86.45 83.883 ;
      RECT 85.748 83.774 86.496 83.837 ;
      RECT 85.794 83.728 86.542 83.791 ;
      RECT 85.84 83.682 86.588 83.745 ;
      RECT 85.886 83.636 86.634 83.699 ;
      RECT 85.932 83.59 86.68 83.653 ;
      RECT 85.978 83.544 86.726 83.607 ;
      RECT 86.024 83.498 86.772 83.561 ;
      RECT 86.07 83.452 86.818 83.515 ;
      RECT 86.116 83.406 86.864 83.469 ;
      RECT 86.162 83.36 86.91 83.423 ;
      RECT 86.208 83.314 86.956 83.377 ;
      RECT 86.254 83.268 87.002 83.331 ;
      RECT 86.3 83.222 87.048 83.285 ;
      RECT 86.346 83.176 87.094 83.239 ;
      RECT 86.392 83.13 87.14 83.193 ;
      RECT 86.438 83.084 87.186 83.147 ;
      RECT 86.484 83.038 87.232 83.101 ;
      RECT 86.53 82.992 87.278 83.055 ;
      RECT 86.576 82.946 87.324 83.009 ;
      RECT 86.622 82.9 87.37 82.963 ;
      RECT 86.668 82.854 87.416 82.917 ;
      RECT 86.714 82.808 87.462 82.871 ;
      RECT 86.76 82.762 87.508 82.825 ;
      RECT 86.806 82.716 87.554 82.779 ;
      RECT 86.852 82.67 87.6 82.733 ;
      RECT 86.898 82.624 87.646 82.687 ;
      RECT 86.944 82.578 87.692 82.641 ;
      RECT 86.99 82.532 87.738 82.595 ;
      RECT 87.036 82.486 87.784 82.549 ;
      RECT 87.082 82.44 87.83 82.503 ;
      RECT 87.128 82.394 87.876 82.457 ;
      RECT 87.174 82.348 87.922 82.411 ;
      RECT 87.22 82.302 87.968 82.365 ;
      RECT 87.266 82.256 88.014 82.319 ;
      RECT 87.312 82.21 88.06 82.273 ;
      RECT 87.358 82.164 88.106 82.227 ;
      RECT 87.404 82.118 88.152 82.181 ;
      RECT 87.45 82.072 88.198 82.135 ;
      RECT 87.496 82.026 88.244 82.089 ;
      RECT 87.542 81.98 88.29 82.043 ;
      RECT 87.588 81.934 88.336 81.997 ;
      RECT 87.634 81.888 88.382 81.951 ;
      RECT 87.68 81.842 88.428 81.905 ;
      RECT 87.726 81.796 88.474 81.859 ;
      RECT 87.772 81.75 88.52 81.813 ;
      RECT 87.818 81.704 88.566 81.767 ;
      RECT 87.864 81.658 88.612 81.721 ;
      RECT 87.91 81.612 88.658 81.675 ;
      RECT 87.956 81.566 88.704 81.629 ;
      RECT 88.692 80.852 88.704 81.629 ;
      RECT 88.002 81.52 88.75 81.583 ;
      RECT 88.695 80.827 88.75 81.583 ;
      RECT 88.048 81.474 88.796 81.537 ;
      RECT 88.741 80.781 88.796 81.537 ;
      RECT 88.094 81.428 88.842 81.491 ;
      RECT 88.787 80.735 88.842 81.491 ;
      RECT 88.14 81.382 88.888 81.445 ;
      RECT 88.833 80.689 88.888 81.445 ;
      RECT 88.186 81.336 88.934 81.399 ;
      RECT 88.879 80.643 88.934 81.399 ;
      RECT 88.232 81.29 88.98 81.353 ;
      RECT 88.925 80.597 88.98 81.353 ;
      RECT 88.278 81.244 89.026 81.307 ;
      RECT 88.971 80.551 89.026 81.307 ;
      RECT 88.324 81.198 89.072 81.261 ;
      RECT 89.017 80.505 89.072 81.261 ;
      RECT 88.37 81.152 89.118 81.215 ;
      RECT 89.063 80.459 89.118 81.215 ;
      RECT 88.416 81.106 89.164 81.169 ;
      RECT 89.109 80.413 89.164 81.169 ;
      RECT 88.416 81.106 89.17 81.143 ;
      RECT 88.462 81.06 89.216 81.117 ;
      RECT 89.155 80.367 89.216 81.117 ;
      RECT 88.508 81.014 89.262 81.071 ;
      RECT 89.201 80.321 89.262 81.071 ;
      RECT 88.554 80.968 89.308 81.025 ;
      RECT 89.247 80.275 89.308 81.025 ;
      RECT 88.6 80.922 89.354 80.979 ;
      RECT 89.293 80.229 89.354 80.979 ;
      RECT 88.646 80.876 89.4 80.933 ;
      RECT 89.339 80.183 89.4 80.933 ;
      RECT 89.385 80.137 89.446 80.887 ;
      RECT 89.431 80.091 89.492 80.841 ;
      RECT 89.477 80.045 89.538 80.795 ;
      RECT 89.523 79.999 89.584 80.749 ;
      RECT 89.569 79.953 89.63 80.703 ;
      RECT 89.615 79.907 89.676 80.657 ;
      RECT 89.661 79.861 89.722 80.611 ;
      RECT 89.707 79.815 89.768 80.565 ;
      RECT 89.753 79.769 89.814 80.519 ;
      RECT 89.799 79.723 89.86 80.473 ;
      RECT 89.845 79.677 89.906 80.427 ;
      RECT 89.891 79.631 89.952 80.381 ;
      RECT 89.937 79.585 89.998 80.335 ;
      RECT 89.983 79.539 90.044 80.289 ;
      RECT 90.029 79.493 90.09 80.243 ;
      RECT 90.075 79.447 90.136 80.197 ;
      RECT 90.121 79.401 90.182 80.151 ;
      RECT 90.167 79.355 90.228 80.105 ;
      RECT 90.213 79.309 90.274 80.059 ;
      RECT 90.259 79.263 90.32 80.013 ;
      RECT 90.305 79.217 90.366 79.967 ;
      RECT 90.351 79.171 90.412 79.921 ;
      RECT 90.397 79.125 90.458 79.875 ;
      RECT 90.443 79.079 90.504 79.829 ;
      RECT 90.489 79.033 90.55 79.783 ;
      RECT 90.535 78.987 90.596 79.737 ;
      RECT 90.581 78.941 90.642 79.691 ;
      RECT 90.627 78.895 90.688 79.645 ;
      RECT 90.673 78.849 90.734 79.599 ;
      RECT 90.719 78.803 90.78 79.553 ;
      RECT 90.765 78.757 90.826 79.507 ;
      RECT 90.811 78.711 90.872 79.461 ;
      RECT 90.857 78.665 90.918 79.415 ;
      RECT 90.903 78.619 90.964 79.369 ;
      RECT 90.949 78.573 91.01 79.323 ;
      RECT 90.995 78.527 91.056 79.277 ;
      RECT 91.041 78.481 91.102 79.231 ;
      RECT 91.087 78.435 91.148 79.185 ;
      RECT 91.133 78.389 91.194 79.139 ;
      RECT 91.179 78.343 91.24 79.093 ;
      RECT 91.225 78.297 91.286 79.047 ;
      RECT 91.271 78.251 91.332 79.001 ;
      RECT 91.317 78.205 91.378 78.955 ;
      RECT 91.363 78.159 91.424 78.909 ;
      RECT 91.409 78.113 91.47 78.863 ;
      RECT 91.455 78.067 91.516 78.817 ;
      RECT 91.501 78.021 91.562 78.771 ;
      RECT 91.547 77.975 91.608 78.725 ;
      RECT 91.593 77.929 91.654 78.679 ;
      RECT 91.639 77.883 91.7 78.633 ;
      RECT 91.685 77.837 91.746 78.587 ;
      RECT 91.731 77.791 91.792 78.541 ;
      RECT 91.777 77.745 91.838 78.495 ;
      RECT 91.823 77.699 91.884 78.449 ;
      RECT 91.869 77.653 91.93 78.403 ;
      RECT 91.915 77.607 91.976 78.357 ;
      RECT 91.961 77.561 92.022 78.311 ;
      RECT 92.007 77.515 92.068 78.265 ;
      RECT 92.053 77.469 92.114 78.219 ;
      RECT 91.363 78.159 92.14 78.183 ;
      RECT 92.215 77.33 110 78.17 ;
      RECT 92.191 77.342 110 78.17 ;
      RECT 92.145 77.377 110 78.17 ;
      RECT 92.099 77.423 110 78.17 ;
      RECT 89.83 97.327 90.67 110 ;
      RECT 89.83 97.327 90.716 99.197 ;
      RECT 89.83 97.327 90.762 99.151 ;
      RECT 89.83 97.327 90.808 99.105 ;
      RECT 89.83 97.327 90.854 99.059 ;
      RECT 89.83 97.327 90.9 99.013 ;
      RECT 89.83 97.327 90.946 98.967 ;
      RECT 89.83 97.327 90.992 98.921 ;
      RECT 89.83 97.327 91.038 98.875 ;
      RECT 89.83 97.327 91.084 98.829 ;
      RECT 89.83 97.327 91.13 98.783 ;
      RECT 89.83 97.327 91.176 98.737 ;
      RECT 89.83 97.327 91.222 98.691 ;
      RECT 89.83 97.327 91.268 98.645 ;
      RECT 89.83 97.327 91.314 98.599 ;
      RECT 89.83 97.327 91.36 98.553 ;
      RECT 89.83 97.327 91.406 98.507 ;
      RECT 89.83 97.327 91.452 98.461 ;
      RECT 89.83 97.327 91.498 98.415 ;
      RECT 89.83 97.327 91.544 98.369 ;
      RECT 89.83 97.327 91.59 98.323 ;
      RECT 89.83 97.327 91.636 98.277 ;
      RECT 89.83 97.327 91.682 98.231 ;
      RECT 89.83 97.327 91.728 98.185 ;
      RECT 89.83 97.327 91.774 98.139 ;
      RECT 89.83 97.327 91.82 98.093 ;
      RECT 89.83 97.327 91.866 98.047 ;
      RECT 89.83 97.327 91.912 98.001 ;
      RECT 89.83 97.327 91.958 97.955 ;
      RECT 89.83 97.327 92.004 97.909 ;
      RECT 89.83 97.327 92.05 97.863 ;
      RECT 89.83 97.327 92.096 97.817 ;
      RECT 89.83 97.327 92.142 97.771 ;
      RECT 89.83 97.327 92.188 97.725 ;
      RECT 89.83 97.327 92.234 97.679 ;
      RECT 89.83 97.327 92.28 97.633 ;
      RECT 89.83 97.327 92.326 97.587 ;
      RECT 89.83 97.327 92.372 97.541 ;
      RECT 89.83 97.327 92.418 97.495 ;
      RECT 89.83 97.327 92.464 97.449 ;
      RECT 89.83 97.327 92.51 97.403 ;
      RECT 89.876 97.281 92.556 97.357 ;
      RECT 92.498 94.659 92.556 97.357 ;
      RECT 89.922 97.235 92.602 97.311 ;
      RECT 92.544 94.613 92.602 97.311 ;
      RECT 89.968 97.189 92.648 97.265 ;
      RECT 92.59 94.567 92.648 97.265 ;
      RECT 90.014 97.143 92.694 97.219 ;
      RECT 92.636 94.521 92.694 97.219 ;
      RECT 90.06 97.097 92.74 97.173 ;
      RECT 92.682 94.475 92.74 97.173 ;
      RECT 90.106 97.051 92.786 97.127 ;
      RECT 92.728 94.429 92.786 97.127 ;
      RECT 90.152 97.005 92.832 97.081 ;
      RECT 92.774 94.393 92.832 97.081 ;
      RECT 90.198 96.959 92.878 97.035 ;
      RECT 92.8 94.357 92.878 97.035 ;
      RECT 90.244 96.913 92.924 96.989 ;
      RECT 92.846 94.311 92.924 96.989 ;
      RECT 90.29 96.867 92.97 96.943 ;
      RECT 92.892 94.265 92.97 96.943 ;
      RECT 90.336 96.821 93.016 96.897 ;
      RECT 92.938 94.219 93.016 96.897 ;
      RECT 90.382 96.775 93.062 96.851 ;
      RECT 92.984 94.173 93.062 96.851 ;
      RECT 90.428 96.729 93.108 96.805 ;
      RECT 93.03 94.127 93.108 96.805 ;
      RECT 90.474 96.683 93.154 96.759 ;
      RECT 93.076 94.081 93.154 96.759 ;
      RECT 90.52 96.637 93.2 96.713 ;
      RECT 93.122 94.035 93.2 96.713 ;
      RECT 90.566 96.591 93.246 96.667 ;
      RECT 93.168 93.989 93.246 96.667 ;
      RECT 90.612 96.545 93.292 96.621 ;
      RECT 93.214 93.943 93.292 96.621 ;
      RECT 90.658 96.499 93.338 96.575 ;
      RECT 93.26 93.897 93.338 96.575 ;
      RECT 90.704 96.453 93.384 96.529 ;
      RECT 93.306 93.851 93.384 96.529 ;
      RECT 90.75 96.407 93.43 96.483 ;
      RECT 93.352 93.805 93.43 96.483 ;
      RECT 90.796 96.361 93.476 96.437 ;
      RECT 93.398 93.759 93.476 96.437 ;
      RECT 90.842 96.315 93.522 96.391 ;
      RECT 93.444 93.713 93.522 96.391 ;
      RECT 90.888 96.269 93.568 96.345 ;
      RECT 93.49 93.667 93.568 96.345 ;
      RECT 90.934 96.223 93.614 96.299 ;
      RECT 93.536 93.621 93.614 96.299 ;
      RECT 90.98 96.177 93.66 96.253 ;
      RECT 93.582 93.575 93.66 96.253 ;
      RECT 91.026 96.131 93.706 96.207 ;
      RECT 93.628 93.529 93.706 96.207 ;
      RECT 91.072 96.085 93.752 96.161 ;
      RECT 93.674 93.483 93.752 96.161 ;
      RECT 91.118 96.039 93.798 96.115 ;
      RECT 93.72 93.437 93.798 96.115 ;
      RECT 91.164 95.993 93.844 96.069 ;
      RECT 93.766 93.391 93.844 96.069 ;
      RECT 91.21 95.947 93.89 96.023 ;
      RECT 93.812 93.345 93.89 96.023 ;
      RECT 91.256 95.901 93.936 95.977 ;
      RECT 93.858 93.299 93.936 95.977 ;
      RECT 91.302 95.855 93.982 95.931 ;
      RECT 93.904 93.253 93.982 95.931 ;
      RECT 91.348 95.809 94.028 95.885 ;
      RECT 93.95 93.207 94.028 95.885 ;
      RECT 91.394 95.763 94.074 95.839 ;
      RECT 93.996 93.161 94.074 95.839 ;
      RECT 91.44 95.717 94.12 95.793 ;
      RECT 94.042 93.115 94.12 95.793 ;
      RECT 91.486 95.671 94.166 95.747 ;
      RECT 94.088 93.069 94.166 95.747 ;
      RECT 91.532 95.625 94.212 95.701 ;
      RECT 94.134 93.023 94.212 95.701 ;
      RECT 91.578 95.579 94.258 95.655 ;
      RECT 94.18 92.977 94.258 95.655 ;
      RECT 91.624 95.533 94.304 95.609 ;
      RECT 94.226 92.931 94.304 95.609 ;
      RECT 91.67 95.487 94.35 95.563 ;
      RECT 94.272 92.885 94.35 95.563 ;
      RECT 91.716 95.441 94.396 95.517 ;
      RECT 94.318 92.839 94.396 95.517 ;
      RECT 91.762 95.395 94.442 95.471 ;
      RECT 94.364 92.793 94.442 95.471 ;
      RECT 91.808 95.349 94.488 95.425 ;
      RECT 94.41 92.747 94.488 95.425 ;
      RECT 91.854 95.303 94.534 95.379 ;
      RECT 94.456 92.701 94.534 95.379 ;
      RECT 91.9 95.257 94.58 95.333 ;
      RECT 94.502 92.655 94.58 95.333 ;
      RECT 91.946 95.211 94.626 95.287 ;
      RECT 94.548 92.609 94.626 95.287 ;
      RECT 91.992 95.165 94.672 95.241 ;
      RECT 94.594 92.563 94.672 95.241 ;
      RECT 92.038 95.119 94.718 95.195 ;
      RECT 94.64 92.517 94.718 95.195 ;
      RECT 92.084 95.073 94.764 95.149 ;
      RECT 94.686 92.471 94.764 95.149 ;
      RECT 92.13 95.027 94.81 95.103 ;
      RECT 94.732 92.425 94.81 95.103 ;
      RECT 92.176 94.981 94.856 95.057 ;
      RECT 94.778 92.379 94.856 95.057 ;
      RECT 92.222 94.935 94.902 95.011 ;
      RECT 94.824 92.333 94.902 95.011 ;
      RECT 92.268 94.889 94.948 94.965 ;
      RECT 94.87 92.287 94.948 94.965 ;
      RECT 92.314 94.843 94.994 94.919 ;
      RECT 94.916 92.241 94.994 94.919 ;
      RECT 92.36 94.797 95.04 94.873 ;
      RECT 94.962 92.195 95.04 94.873 ;
      RECT 92.406 94.751 95.086 94.827 ;
      RECT 95.008 92.149 95.086 94.827 ;
      RECT 92.452 94.705 95.132 94.781 ;
      RECT 95.054 92.103 95.132 94.781 ;
      RECT 95.1 92.057 95.178 94.735 ;
      RECT 95.146 92.011 95.224 94.689 ;
      RECT 95.192 91.965 95.27 94.643 ;
      RECT 95.238 91.919 95.316 94.597 ;
      RECT 95.284 91.873 95.362 94.551 ;
      RECT 95.33 91.827 95.408 94.505 ;
      RECT 95.376 91.781 95.454 94.459 ;
      RECT 95.422 91.735 95.5 94.413 ;
      RECT 95.468 91.689 95.546 94.367 ;
      RECT 95.514 91.643 95.592 94.321 ;
      RECT 95.56 91.597 95.638 94.275 ;
      RECT 95.606 91.551 95.684 94.229 ;
      RECT 95.652 91.505 95.73 94.183 ;
      RECT 95.698 91.459 95.776 94.137 ;
      RECT 95.744 91.413 95.822 94.091 ;
      RECT 95.79 91.367 95.868 94.045 ;
      RECT 95.836 91.321 95.914 93.999 ;
      RECT 95.882 91.275 95.96 93.953 ;
      RECT 95.928 91.229 96.006 93.907 ;
      RECT 95.974 91.183 96.052 93.861 ;
      RECT 96.02 91.137 96.098 93.815 ;
      RECT 96.066 91.091 96.144 93.769 ;
      RECT 96.112 91.045 96.19 93.723 ;
      RECT 96.158 90.999 96.236 93.677 ;
      RECT 96.204 90.953 96.282 93.631 ;
      RECT 96.25 90.907 96.328 93.585 ;
      RECT 96.296 90.861 96.374 93.539 ;
      RECT 96.342 90.815 96.42 93.493 ;
      RECT 96.388 90.769 96.466 93.447 ;
      RECT 96.434 90.723 96.512 93.401 ;
      RECT 96.48 90.677 96.558 93.355 ;
      RECT 96.526 90.631 96.604 93.309 ;
      RECT 96.572 90.585 96.65 93.263 ;
      RECT 96.618 90.539 96.696 93.217 ;
      RECT 96.664 90.493 96.742 93.171 ;
      RECT 96.71 90.447 96.788 93.125 ;
      RECT 96.756 90.401 96.834 93.079 ;
      RECT 96.802 90.355 96.88 93.033 ;
      RECT 96.848 90.309 96.926 92.987 ;
      RECT 96.894 90.263 96.972 92.941 ;
      RECT 96.94 90.217 97.018 92.895 ;
      RECT 96.986 90.171 97.064 92.849 ;
      RECT 97.032 90.125 97.11 92.803 ;
      RECT 97.078 90.079 97.156 92.757 ;
      RECT 97.124 90.033 97.202 92.711 ;
      RECT 97.17 89.987 97.248 92.665 ;
      RECT 97.216 89.941 97.294 92.619 ;
      RECT 97.262 89.895 97.34 92.573 ;
      RECT 97.308 89.851 97.386 92.527 ;
      RECT 97.35 89.83 97.432 92.481 ;
      RECT 97.35 89.83 97.478 92.435 ;
      RECT 97.35 89.83 97.524 92.389 ;
      RECT 97.35 89.83 97.57 92.343 ;
      RECT 97.35 89.83 97.616 92.297 ;
      RECT 97.35 89.83 97.662 92.251 ;
      RECT 94.962 92.195 97.67 92.224 ;
      RECT 97.35 89.83 97.716 92.197 ;
      RECT 97.35 89.83 97.762 92.151 ;
      RECT 97.35 89.83 97.808 92.105 ;
      RECT 97.35 89.83 97.854 92.059 ;
      RECT 97.35 89.83 97.9 92.013 ;
      RECT 97.35 89.83 97.946 91.967 ;
      RECT 97.35 89.83 97.992 91.921 ;
      RECT 97.35 89.83 98.038 91.875 ;
      RECT 97.35 89.83 98.084 91.829 ;
      RECT 97.35 89.83 98.13 91.783 ;
      RECT 97.35 89.83 98.176 91.737 ;
      RECT 97.35 89.83 98.222 91.691 ;
      RECT 97.35 89.83 98.268 91.645 ;
      RECT 97.35 89.83 98.314 91.599 ;
      RECT 97.35 89.83 98.36 91.553 ;
      RECT 97.35 89.83 98.406 91.507 ;
      RECT 97.35 89.83 98.452 91.461 ;
      RECT 97.35 89.83 98.498 91.415 ;
      RECT 97.35 89.83 98.544 91.369 ;
      RECT 97.35 89.83 98.59 91.323 ;
      RECT 97.35 89.83 98.636 91.277 ;
      RECT 97.35 89.83 98.682 91.231 ;
      RECT 97.35 89.83 98.728 91.185 ;
      RECT 97.35 89.83 98.774 91.139 ;
      RECT 97.35 89.83 98.82 91.093 ;
      RECT 97.35 89.83 98.866 91.047 ;
      RECT 97.35 89.83 98.912 91.001 ;
      RECT 97.35 89.83 98.958 90.955 ;
      RECT 97.35 89.83 99.004 90.909 ;
      RECT 97.35 89.83 99.05 90.863 ;
      RECT 97.35 89.83 99.096 90.817 ;
      RECT 97.35 89.83 99.142 90.771 ;
      RECT 97.35 89.83 99.188 90.725 ;
      RECT 97.35 89.83 99.22 90.686 ;
      RECT 97.35 89.83 110 90.67 ;
      RECT 98.33 102.757 99.17 110 ;
      RECT 98.33 102.757 99.216 103.487 ;
      RECT 98.33 102.757 99.262 103.441 ;
      RECT 98.33 102.757 99.308 103.395 ;
      RECT 98.33 102.757 99.354 103.349 ;
      RECT 98.33 102.757 99.4 103.303 ;
      RECT 98.33 102.757 99.446 103.257 ;
      RECT 98.33 102.757 99.492 103.211 ;
      RECT 98.33 102.757 99.538 103.165 ;
      RECT 98.33 102.757 99.584 103.119 ;
      RECT 98.33 102.757 99.63 103.073 ;
      RECT 98.33 102.757 99.676 103.027 ;
      RECT 98.33 102.757 99.722 102.981 ;
      RECT 98.33 102.757 99.768 102.935 ;
      RECT 98.33 102.757 99.814 102.889 ;
      RECT 98.33 102.757 99.86 102.843 ;
      RECT 98.376 102.711 99.906 102.797 ;
      RECT 99.848 101.246 99.906 102.797 ;
      RECT 98.422 102.665 99.952 102.751 ;
      RECT 99.88 101.207 99.952 102.751 ;
      RECT 98.468 102.619 99.998 102.705 ;
      RECT 99.926 101.161 99.998 102.705 ;
      RECT 98.514 102.573 100.044 102.659 ;
      RECT 99.972 101.115 100.044 102.659 ;
      RECT 98.56 102.527 100.09 102.613 ;
      RECT 100.018 101.069 100.09 102.613 ;
      RECT 98.606 102.481 100.136 102.567 ;
      RECT 100.064 101.023 100.136 102.567 ;
      RECT 98.652 102.435 100.182 102.521 ;
      RECT 100.11 100.977 100.182 102.521 ;
      RECT 98.698 102.389 100.228 102.475 ;
      RECT 100.156 100.931 100.228 102.475 ;
      RECT 98.744 102.343 100.274 102.429 ;
      RECT 100.202 100.885 100.274 102.429 ;
      RECT 98.79 102.297 100.32 102.383 ;
      RECT 100.248 100.839 100.32 102.383 ;
      RECT 98.836 102.251 100.366 102.337 ;
      RECT 100.294 100.793 100.366 102.337 ;
      RECT 98.882 102.205 100.412 102.291 ;
      RECT 100.34 100.747 100.412 102.291 ;
      RECT 98.928 102.159 100.458 102.245 ;
      RECT 100.386 100.701 100.458 102.245 ;
      RECT 98.974 102.113 100.504 102.199 ;
      RECT 100.432 100.655 100.504 102.199 ;
      RECT 99.02 102.067 100.55 102.153 ;
      RECT 100.478 100.609 100.55 102.153 ;
      RECT 99.066 102.021 100.596 102.107 ;
      RECT 100.524 100.563 100.596 102.107 ;
      RECT 99.112 101.975 100.642 102.061 ;
      RECT 100.57 100.517 100.642 102.061 ;
      RECT 99.158 101.929 100.688 102.015 ;
      RECT 100.616 100.471 100.688 102.015 ;
      RECT 99.204 101.883 100.734 101.969 ;
      RECT 100.662 100.425 100.734 101.969 ;
      RECT 99.25 101.837 100.78 101.923 ;
      RECT 100.708 100.379 100.78 101.923 ;
      RECT 99.296 101.791 100.826 101.877 ;
      RECT 100.754 100.333 100.826 101.877 ;
      RECT 99.342 101.745 100.872 101.831 ;
      RECT 100.8 100.287 100.872 101.831 ;
      RECT 99.388 101.699 100.918 101.785 ;
      RECT 100.846 100.241 100.918 101.785 ;
      RECT 99.434 101.653 100.964 101.739 ;
      RECT 100.892 100.195 100.964 101.739 ;
      RECT 99.48 101.607 101.01 101.693 ;
      RECT 100.938 100.149 101.01 101.693 ;
      RECT 99.526 101.561 101.056 101.647 ;
      RECT 100.984 100.103 101.056 101.647 ;
      RECT 99.572 101.515 101.102 101.601 ;
      RECT 101.03 100.057 101.102 101.601 ;
      RECT 99.618 101.469 101.148 101.555 ;
      RECT 101.076 100.011 101.148 101.555 ;
      RECT 99.664 101.423 101.194 101.509 ;
      RECT 101.122 99.965 101.194 101.509 ;
      RECT 99.71 101.377 101.24 101.463 ;
      RECT 101.168 99.919 101.24 101.463 ;
      RECT 99.756 101.331 101.286 101.417 ;
      RECT 101.214 99.873 101.286 101.417 ;
      RECT 99.802 101.285 101.332 101.371 ;
      RECT 101.26 99.827 101.332 101.371 ;
      RECT 101.306 99.781 101.378 101.325 ;
      RECT 101.352 99.735 101.424 101.279 ;
      RECT 101.398 99.689 101.47 101.233 ;
      RECT 101.444 99.643 101.516 101.187 ;
      RECT 101.49 99.597 101.562 101.141 ;
      RECT 101.536 99.551 101.608 101.095 ;
      RECT 101.582 99.505 101.654 101.049 ;
      RECT 101.628 99.459 101.7 101.003 ;
      RECT 101.674 99.413 101.746 100.957 ;
      RECT 101.72 99.367 101.792 100.911 ;
      RECT 101.766 99.321 101.838 100.865 ;
      RECT 101.812 99.275 101.884 100.819 ;
      RECT 101.858 99.229 101.93 100.773 ;
      RECT 101.904 99.183 101.976 100.727 ;
      RECT 101.95 99.137 102.022 100.681 ;
      RECT 101.996 99.091 102.068 100.635 ;
      RECT 102.042 99.045 102.114 100.589 ;
      RECT 102.088 98.999 102.16 100.543 ;
      RECT 102.134 98.953 102.206 100.497 ;
      RECT 102.18 98.907 102.252 100.451 ;
      RECT 102.226 98.861 102.298 100.405 ;
      RECT 102.272 98.815 102.344 100.359 ;
      RECT 102.318 98.769 102.39 100.313 ;
      RECT 102.364 98.723 102.436 100.267 ;
      RECT 102.41 98.677 102.482 100.221 ;
      RECT 102.456 98.631 102.528 100.175 ;
      RECT 102.502 98.585 102.574 100.129 ;
      RECT 102.548 98.539 102.62 100.083 ;
      RECT 102.594 98.493 102.666 100.037 ;
      RECT 102.64 98.447 102.712 99.991 ;
      RECT 102.686 98.401 102.758 99.945 ;
      RECT 102.732 98.354 102.804 99.899 ;
      RECT 102.778 98.33 102.85 99.853 ;
      RECT 102.778 98.33 102.896 99.807 ;
      RECT 102.778 98.33 102.942 99.761 ;
      RECT 102.778 98.33 102.988 99.715 ;
      RECT 102.778 98.33 103.034 99.669 ;
      RECT 102.778 98.33 103.08 99.623 ;
      RECT 102.778 98.33 103.126 99.577 ;
      RECT 102.778 98.33 103.172 99.531 ;
      RECT 102.778 98.33 103.218 99.485 ;
      RECT 102.778 98.33 103.264 99.439 ;
      RECT 102.778 98.33 103.31 99.393 ;
      RECT 102.778 98.33 103.356 99.347 ;
      RECT 102.778 98.33 103.402 99.301 ;
      RECT 102.778 98.33 103.448 99.255 ;
      RECT 102.778 98.33 103.494 99.209 ;
      RECT 101.95 99.137 103.51 99.178 ;
      RECT 102.778 98.33 110 99.17 ;
      RECT 107.83 109.057 110 110 ;
      RECT 109.08 107.83 110 110 ;
      RECT 107.876 109.011 110 110 ;
      RECT 109.072 107.834 110 110 ;
      RECT 107.922 108.965 110 110 ;
      RECT 109.026 107.861 110 110 ;
      RECT 107.968 108.919 110 110 ;
      RECT 108.98 107.907 110 110 ;
      RECT 108.014 108.873 110 110 ;
      RECT 108.934 107.953 110 110 ;
      RECT 108.06 108.827 110 110 ;
      RECT 108.888 107.999 110 110 ;
      RECT 108.106 108.781 110 110 ;
      RECT 108.842 108.045 110 110 ;
      RECT 108.152 108.735 110 110 ;
      RECT 108.796 108.091 110 110 ;
      RECT 108.198 108.689 110 110 ;
      RECT 108.75 108.137 110 110 ;
      RECT 108.244 108.643 110 110 ;
      RECT 108.704 108.183 110 110 ;
      RECT 108.29 108.597 110 110 ;
      RECT 108.658 108.229 110 110 ;
      RECT 108.336 108.551 110 110 ;
      RECT 108.612 108.275 110 110 ;
      RECT 108.382 108.505 110 110 ;
      RECT 108.566 108.321 110 110 ;
      RECT 108.428 108.459 110 110 ;
      RECT 108.52 108.367 110 110 ;
      RECT 108.474 108.413 110 110 ;
    LAYER T4M2 SPACING 0.4 ;
      RECT -20 -20 2.9 110 ;
      RECT -20 -20 2.946 55.392 ;
      RECT -20 -20 2.992 55.346 ;
      RECT -20 -20 3.038 55.3 ;
      RECT -20 -20 3.084 55.254 ;
      RECT -20 -20 3.13 55.208 ;
      RECT -20 -20 3.176 55.162 ;
      RECT -20 -20 3.222 55.116 ;
      RECT -20 -20 3.268 55.07 ;
      RECT -20 -20 3.314 55.024 ;
      RECT -20 -20 3.36 54.978 ;
      RECT -20 -20 3.406 54.932 ;
      RECT -20 -20 3.452 54.886 ;
      RECT -20 -20 3.498 54.84 ;
      RECT -20 -20 3.544 54.794 ;
      RECT -20 -20 3.59 54.748 ;
      RECT -20 -20 3.636 54.702 ;
      RECT -20 -20 3.682 54.656 ;
      RECT -20 -20 3.728 54.61 ;
      RECT -20 -20 3.774 54.564 ;
      RECT -20 -20 3.82 54.518 ;
      RECT -20 -20 3.866 54.472 ;
      RECT -20 -20 3.912 54.426 ;
      RECT -20 -20 3.958 54.38 ;
      RECT -20 -20 4.004 54.334 ;
      RECT -20 -20 4.05 54.288 ;
      RECT -20 -20 4.096 54.242 ;
      RECT -20 -20 4.142 54.196 ;
      RECT -20 -20 4.188 54.15 ;
      RECT -20 -20 4.234 54.104 ;
      RECT -20 -20 4.28 54.058 ;
      RECT -20 -20 4.326 54.012 ;
      RECT -20 -20 4.372 53.966 ;
      RECT -20 -20 4.418 53.92 ;
      RECT -20 -20 4.464 53.874 ;
      RECT -20 -20 4.51 53.828 ;
      RECT -20 -20 4.556 53.782 ;
      RECT -20 -20 4.602 53.736 ;
      RECT -20 -20 4.648 53.69 ;
      RECT -20 -20 4.694 53.644 ;
      RECT -20 -20 4.74 53.598 ;
      RECT -20 -20 4.786 53.552 ;
      RECT -20 -20 4.832 53.506 ;
      RECT -20 -20 4.878 53.46 ;
      RECT -20 -20 4.924 53.414 ;
      RECT -20 -20 4.97 53.368 ;
      RECT -20 -20 5.016 53.322 ;
      RECT -20 -20 5.062 53.276 ;
      RECT -20 -20 5.108 53.23 ;
      RECT -20 -20 5.154 53.184 ;
      RECT -20 -20 5.2 53.138 ;
      RECT -20 -20 5.246 53.092 ;
      RECT -20 -20 5.292 53.046 ;
      RECT -20 -20 5.338 53 ;
      RECT -20 -20 5.384 52.954 ;
      RECT -20 -20 5.43 52.908 ;
      RECT -20 -20 5.476 52.862 ;
      RECT -20 -20 5.522 52.816 ;
      RECT -20 -20 5.568 52.77 ;
      RECT -20 -20 5.614 52.724 ;
      RECT -20 -20 5.66 52.678 ;
      RECT -20 -20 5.706 52.632 ;
      RECT -20 -20 5.752 52.586 ;
      RECT -20 -20 5.798 52.54 ;
      RECT -20 -20 5.844 52.494 ;
      RECT -20 -20 5.89 52.448 ;
      RECT -20 -20 5.936 52.402 ;
      RECT -20 -20 5.982 52.356 ;
      RECT -20 -20 6.028 52.31 ;
      RECT -20 -20 6.074 52.264 ;
      RECT -20 -20 6.12 52.218 ;
      RECT -20 -20 6.166 52.172 ;
      RECT -20 -20 6.212 52.126 ;
      RECT -20 -20 6.258 52.08 ;
      RECT -20 -20 6.304 52.034 ;
      RECT -20 -20 6.35 51.988 ;
      RECT -20 -20 6.396 51.942 ;
      RECT -20 -20 6.442 51.896 ;
      RECT -20 -20 6.488 51.85 ;
      RECT -20 -20 6.534 51.804 ;
      RECT -20 -20 6.58 51.758 ;
      RECT -20 -20 6.626 51.712 ;
      RECT -20 -20 6.672 51.666 ;
      RECT -20 -20 6.718 51.62 ;
      RECT -20 -20 6.764 51.574 ;
      RECT -20 -20 6.81 51.528 ;
      RECT -20 -20 6.856 51.482 ;
      RECT -20 -20 6.902 51.436 ;
      RECT -20 -20 6.948 51.39 ;
      RECT -20 -20 6.994 51.344 ;
      RECT -20 -20 7.04 51.298 ;
      RECT -20 -20 7.086 51.252 ;
      RECT -20 -20 7.132 51.206 ;
      RECT -20 -20 7.178 51.16 ;
      RECT -20 -20 7.224 51.114 ;
      RECT -20 -20 7.27 51.068 ;
      RECT -20 -20 7.316 51.022 ;
      RECT -20 -20 7.362 50.976 ;
      RECT -20 -20 7.408 50.93 ;
      RECT -20 -20 7.454 50.884 ;
      RECT -20 -20 7.5 50.838 ;
      RECT -20 -20 7.546 50.792 ;
      RECT -20 -20 7.592 50.746 ;
      RECT -20 -20 7.638 50.7 ;
      RECT -20 -20 7.684 50.654 ;
      RECT -20 -20 7.73 50.608 ;
      RECT -20 -20 7.776 50.562 ;
      RECT -20 -20 7.822 50.516 ;
      RECT -20 -20 7.868 50.47 ;
      RECT -20 -20 7.914 50.424 ;
      RECT -20 -20 7.96 50.378 ;
      RECT -20 -20 8.006 50.332 ;
      RECT -20 -20 8.052 50.286 ;
      RECT -20 -20 8.098 50.24 ;
      RECT -20 -20 8.144 50.194 ;
      RECT -20 -20 8.19 50.148 ;
      RECT -20 -20 8.236 50.102 ;
      RECT -20 -20 8.282 50.056 ;
      RECT -20 -20 8.328 50.01 ;
      RECT -20 -20 8.374 49.964 ;
      RECT -20 -20 8.42 49.918 ;
      RECT -20 -20 8.466 49.872 ;
      RECT -20 -20 8.512 49.826 ;
      RECT -20 -20 8.558 49.78 ;
      RECT -20 -20 8.604 49.734 ;
      RECT -20 -20 8.65 49.688 ;
      RECT -20 -20 8.696 49.642 ;
      RECT -20 -20 8.742 49.596 ;
      RECT -20 -20 8.788 49.55 ;
      RECT -20 -20 8.834 49.504 ;
      RECT -20 -20 8.88 49.458 ;
      RECT -20 -20 8.926 49.412 ;
      RECT -20 -20 8.972 49.366 ;
      RECT -20 -20 9.018 49.32 ;
      RECT -20 -20 9.064 49.274 ;
      RECT -20 -20 9.11 49.228 ;
      RECT -20 -20 9.156 49.182 ;
      RECT -20 -20 9.202 49.136 ;
      RECT -20 -20 9.248 49.09 ;
      RECT -20 -20 9.294 49.044 ;
      RECT -20 -20 9.34 48.998 ;
      RECT -20 -20 9.386 48.952 ;
      RECT -20 -20 9.432 48.906 ;
      RECT -20 -20 9.478 48.86 ;
      RECT -20 -20 9.524 48.814 ;
      RECT -20 -20 9.57 48.768 ;
      RECT -20 -20 9.616 48.722 ;
      RECT -20 -20 9.662 48.676 ;
      RECT -20 -20 9.708 48.63 ;
      RECT -20 -20 9.754 48.584 ;
      RECT -20 -20 9.8 48.538 ;
      RECT -20 -20 9.846 48.492 ;
      RECT -20 -20 9.892 48.446 ;
      RECT -20 -20 9.938 48.4 ;
      RECT -20 -20 9.984 48.354 ;
      RECT -20 -20 10.03 48.308 ;
      RECT -20 -20 10.076 48.262 ;
      RECT -20 -20 10.122 48.216 ;
      RECT -20 -20 10.168 48.17 ;
      RECT -20 -20 10.214 48.124 ;
      RECT -20 -20 10.26 48.078 ;
      RECT -20 -20 10.306 48.032 ;
      RECT -20 -20 10.352 47.986 ;
      RECT -20 -20 10.398 47.94 ;
      RECT -20 -20 10.444 47.894 ;
      RECT -20 -20 10.49 47.848 ;
      RECT -20 -20 10.536 47.802 ;
      RECT -20 -20 10.582 47.756 ;
      RECT -20 -20 10.628 47.71 ;
      RECT -20 -20 10.674 47.664 ;
      RECT -20 -20 10.72 47.618 ;
      RECT -20 -20 10.766 47.572 ;
      RECT -20 -20 10.812 47.526 ;
      RECT -20 -20 10.858 47.48 ;
      RECT -20 -20 10.904 47.434 ;
      RECT -20 -20 10.95 47.388 ;
      RECT -20 -20 10.996 47.342 ;
      RECT -20 -20 11.042 47.296 ;
      RECT -20 -20 11.088 47.25 ;
      RECT -20 -20 11.134 47.204 ;
      RECT -20 -20 11.18 47.158 ;
      RECT -20 -20 11.226 47.112 ;
      RECT -20 -20 11.272 47.066 ;
      RECT -20 -20 11.318 47.02 ;
      RECT -20 -20 11.364 46.974 ;
      RECT -20 -20 11.41 46.928 ;
      RECT -20 -20 11.456 46.882 ;
      RECT -20 -20 11.502 46.836 ;
      RECT -20 -20 11.548 46.79 ;
      RECT -20 -20 11.594 46.744 ;
      RECT -20 -20 11.64 46.698 ;
      RECT -20 -20 11.686 46.652 ;
      RECT -20 -20 11.732 46.606 ;
      RECT -20 -20 11.778 46.56 ;
      RECT -20 -20 11.824 46.514 ;
      RECT -20 -20 11.87 46.468 ;
      RECT -20 -20 11.916 46.422 ;
      RECT -20 -20 11.962 46.376 ;
      RECT -20 -20 12.008 46.33 ;
      RECT -20 -20 12.054 46.284 ;
      RECT -20 -20 12.1 46.238 ;
      RECT -20 -20 12.146 46.192 ;
      RECT -20 -20 12.192 46.146 ;
      RECT -20 -20 12.238 46.1 ;
      RECT -20 -20 12.284 46.054 ;
      RECT -20 -20 12.33 46.008 ;
      RECT -20 -20 12.376 45.962 ;
      RECT -20 -20 12.422 45.916 ;
      RECT -20 -20 12.468 45.87 ;
      RECT -20 -20 12.514 45.824 ;
      RECT -20 -20 12.56 45.778 ;
      RECT -20 -20 12.606 45.732 ;
      RECT -20 -20 12.652 45.686 ;
      RECT -20 -20 12.698 45.64 ;
      RECT -20 -20 12.744 45.594 ;
      RECT -20 -20 12.79 45.548 ;
      RECT -20 -20 12.836 45.502 ;
      RECT -20 -20 12.882 45.456 ;
      RECT -20 -20 12.928 45.41 ;
      RECT -20 -20 12.974 45.364 ;
      RECT -20 -20 13.02 45.318 ;
      RECT -20 -20 13.066 45.272 ;
      RECT -20 -20 13.112 45.226 ;
      RECT -20 -20 13.158 45.18 ;
      RECT -20 -20 13.204 45.134 ;
      RECT -20 -20 13.25 45.088 ;
      RECT -20 -20 13.296 45.042 ;
      RECT -20 -20 13.342 44.996 ;
      RECT -20 -20 13.388 44.95 ;
      RECT -20 -20 13.434 44.904 ;
      RECT -20 -20 13.48 44.858 ;
      RECT -20 -20 13.526 44.812 ;
      RECT -20 -20 13.572 44.766 ;
      RECT -20 -20 13.618 44.72 ;
      RECT -20 -20 13.664 44.674 ;
      RECT -20 -20 13.71 44.628 ;
      RECT -20 -20 13.756 44.582 ;
      RECT -20 -20 13.802 44.536 ;
      RECT -20 -20 13.848 44.49 ;
      RECT -20 -20 13.894 44.444 ;
      RECT -20 -20 13.94 44.398 ;
      RECT -20 -20 13.986 44.352 ;
      RECT -20 -20 14.032 44.306 ;
      RECT -20 -20 14.078 44.26 ;
      RECT -20 -20 14.124 44.214 ;
      RECT -20 -20 14.17 44.168 ;
      RECT -20 -20 14.216 44.122 ;
      RECT -20 -20 14.262 44.076 ;
      RECT -20 -20 14.308 44.03 ;
      RECT -20 -20 14.354 43.984 ;
      RECT -20 -20 14.4 43.938 ;
      RECT -20 -20 14.446 43.892 ;
      RECT -20 -20 14.492 43.846 ;
      RECT -20 -20 14.538 43.8 ;
      RECT -20 -20 14.584 43.754 ;
      RECT -20 -20 14.63 43.708 ;
      RECT -20 -20 14.676 43.662 ;
      RECT -20 -20 14.722 43.616 ;
      RECT -20 -20 14.768 43.57 ;
      RECT -20 -20 14.814 43.524 ;
      RECT -20 -20 14.86 43.478 ;
      RECT -20 -20 14.9 43.435 ;
      RECT -20 -20 14.946 43.392 ;
      RECT -20 -20 14.992 43.346 ;
      RECT -20 -20 15.038 43.3 ;
      RECT -20 -20 15.084 43.254 ;
      RECT -20 -20 15.13 43.208 ;
      RECT -20 -20 15.176 43.162 ;
      RECT -20 -20 15.222 43.116 ;
      RECT -20 -20 15.268 43.07 ;
      RECT -20 -20 15.314 43.024 ;
      RECT -20 -20 15.36 42.978 ;
      RECT -20 -20 15.406 42.932 ;
      RECT -20 -20 15.452 42.886 ;
      RECT -20 -20 15.498 42.84 ;
      RECT -20 -20 15.544 42.794 ;
      RECT -20 -20 15.59 42.748 ;
      RECT -20 -20 15.636 42.702 ;
      RECT -20 -20 15.682 42.656 ;
      RECT -20 -20 15.728 42.61 ;
      RECT -20 -20 15.774 42.564 ;
      RECT -20 -20 15.82 42.518 ;
      RECT -20 -20 15.866 42.472 ;
      RECT -20 -20 15.912 42.426 ;
      RECT -20 -20 15.958 42.38 ;
      RECT -20 -20 16.004 42.334 ;
      RECT -20 -20 16.05 42.288 ;
      RECT -20 -20 16.096 42.242 ;
      RECT -20 -20 16.142 42.196 ;
      RECT -20 -20 16.188 42.15 ;
      RECT -20 -20 16.234 42.104 ;
      RECT -20 -20 16.28 42.058 ;
      RECT -20 -20 16.326 42.012 ;
      RECT -20 -20 16.372 41.966 ;
      RECT -20 -20 16.418 41.92 ;
      RECT -20 -20 16.464 41.874 ;
      RECT -20 -20 16.51 41.828 ;
      RECT -20 -20 16.556 41.782 ;
      RECT -20 -20 16.602 41.736 ;
      RECT -20 -20 16.648 41.69 ;
      RECT -20 -20 16.694 41.644 ;
      RECT -20 -20 16.74 41.598 ;
      RECT -20 -20 16.786 41.552 ;
      RECT -20 -20 16.832 41.506 ;
      RECT -20 -20 16.878 41.46 ;
      RECT -20 -20 16.924 41.414 ;
      RECT -20 -20 16.97 41.368 ;
      RECT -20 -20 17.016 41.322 ;
      RECT -20 -20 17.062 41.276 ;
      RECT -20 -20 17.108 41.23 ;
      RECT -20 -20 17.154 41.184 ;
      RECT -20 -20 17.2 41.138 ;
      RECT -20 -20 17.246 41.092 ;
      RECT -20 -20 17.292 41.046 ;
      RECT -20 -20 17.338 41 ;
      RECT -20 -20 17.384 40.954 ;
      RECT -20 -20 17.43 40.908 ;
      RECT -20 -20 17.476 40.862 ;
      RECT -20 -20 17.522 40.816 ;
      RECT -20 -20 17.568 40.77 ;
      RECT -20 -20 17.614 40.724 ;
      RECT -20 -20 17.66 40.678 ;
      RECT -20 -20 17.706 40.632 ;
      RECT -20 -20 17.752 40.586 ;
      RECT -20 -20 17.798 40.54 ;
      RECT -20 -20 17.844 40.494 ;
      RECT -20 -20 17.89 40.448 ;
      RECT -20 -20 17.936 40.402 ;
      RECT -20 -20 17.982 40.356 ;
      RECT -20 -20 18.028 40.31 ;
      RECT -20 -20 18.074 40.264 ;
      RECT -20 -20 18.12 40.218 ;
      RECT -20 -20 18.166 40.172 ;
      RECT -20 -20 18.212 40.126 ;
      RECT -20 -20 18.258 40.08 ;
      RECT -20 -20 18.304 40.034 ;
      RECT -20 -20 18.35 39.988 ;
      RECT -20 -20 18.396 39.942 ;
      RECT -20 -20 18.442 39.896 ;
      RECT -20 -20 18.488 39.85 ;
      RECT -20 -20 18.534 39.804 ;
      RECT -20 -20 18.58 39.758 ;
      RECT -20 -20 18.626 39.712 ;
      RECT -20 -20 18.672 39.666 ;
      RECT -20 -20 18.718 39.62 ;
      RECT -20 -20 18.764 39.574 ;
      RECT -20 -20 18.81 39.528 ;
      RECT -20 -20 18.856 39.482 ;
      RECT -20 -20 18.902 39.436 ;
      RECT -20 -20 18.948 39.39 ;
      RECT -20 -20 18.994 39.344 ;
      RECT -20 -20 19.04 39.298 ;
      RECT -20 -20 19.086 39.252 ;
      RECT -20 -20 19.132 39.206 ;
      RECT -20 -20 19.178 39.16 ;
      RECT -20 -20 19.224 39.114 ;
      RECT -20 -20 19.27 39.068 ;
      RECT -20 -20 19.316 39.022 ;
      RECT -20 -20 19.362 38.976 ;
      RECT -20 -20 19.408 38.93 ;
      RECT -20 -20 19.454 38.884 ;
      RECT -20 -20 19.5 38.838 ;
      RECT -20 -20 19.546 38.792 ;
      RECT -20 -20 19.592 38.746 ;
      RECT -20 -20 19.638 38.7 ;
      RECT -20 -20 19.684 38.654 ;
      RECT -20 -20 19.73 38.608 ;
      RECT -20 -20 19.776 38.562 ;
      RECT -20 -20 19.822 38.516 ;
      RECT -20 -20 19.868 38.47 ;
      RECT -20 -20 19.914 38.424 ;
      RECT -20 -20 19.96 38.378 ;
      RECT -20 -20 20.006 38.332 ;
      RECT -20 -20 20.052 38.286 ;
      RECT -20 -20 20.098 38.24 ;
      RECT -20 -20 20.144 38.194 ;
      RECT -20 -20 20.19 38.148 ;
      RECT -20 -20 20.236 38.102 ;
      RECT -20 -20 20.282 38.056 ;
      RECT -20 -20 20.328 38.01 ;
      RECT -20 -20 20.374 37.964 ;
      RECT -20 -20 20.42 37.918 ;
      RECT -20 -20 20.466 37.872 ;
      RECT -20 -20 20.512 37.826 ;
      RECT -20 -20 20.558 37.78 ;
      RECT -20 -20 20.604 37.734 ;
      RECT -20 -20 20.65 37.688 ;
      RECT -20 -20 20.696 37.642 ;
      RECT -20 -20 20.742 37.596 ;
      RECT -20 -20 20.788 37.55 ;
      RECT -20 -20 20.834 37.504 ;
      RECT -20 -20 20.88 37.458 ;
      RECT -20 -20 20.926 37.412 ;
      RECT -20 -20 20.972 37.366 ;
      RECT -20 -20 21.018 37.32 ;
      RECT -20 -20 21.064 37.274 ;
      RECT -20 -20 21.11 37.228 ;
      RECT -20 -20 21.156 37.182 ;
      RECT -20 -20 21.202 37.136 ;
      RECT -20 -20 21.248 37.09 ;
      RECT -20 -20 21.294 37.044 ;
      RECT -20 -20 21.34 36.998 ;
      RECT -20 -20 21.386 36.952 ;
      RECT -20 -20 21.432 36.906 ;
      RECT -20 -20 21.478 36.86 ;
      RECT -20 -20 21.524 36.814 ;
      RECT -20 -20 21.57 36.768 ;
      RECT -20 -20 21.616 36.722 ;
      RECT -20 -20 21.662 36.676 ;
      RECT -20 -20 21.708 36.63 ;
      RECT -20 -20 21.754 36.584 ;
      RECT -20 -20 21.8 36.538 ;
      RECT -20 -20 21.846 36.492 ;
      RECT -20 -20 21.892 36.446 ;
      RECT -20 -20 21.938 36.4 ;
      RECT -20 -20 21.984 36.354 ;
      RECT -20 -20 22.03 36.308 ;
      RECT -20 -20 22.076 36.262 ;
      RECT -20 -20 22.122 36.216 ;
      RECT -20 -20 22.168 36.17 ;
      RECT -20 -20 22.214 36.124 ;
      RECT -20 -20 22.26 36.078 ;
      RECT -20 -20 22.306 36.032 ;
      RECT -20 -20 22.352 35.986 ;
      RECT -20 -20 22.398 35.94 ;
      RECT -20 -20 22.444 35.894 ;
      RECT -20 -20 22.49 35.848 ;
      RECT -20 -20 22.536 35.802 ;
      RECT -20 -20 22.582 35.756 ;
      RECT -20 -20 22.628 35.71 ;
      RECT -20 -20 22.674 35.664 ;
      RECT -20 -20 22.72 35.618 ;
      RECT -20 -20 22.766 35.572 ;
      RECT -20 -20 22.812 35.526 ;
      RECT -20 -20 22.858 35.48 ;
      RECT -20 -20 22.904 35.434 ;
      RECT -20 -20 22.95 35.388 ;
      RECT -20 -20 22.996 35.342 ;
      RECT -20 -20 23.042 35.296 ;
      RECT -20 -20 23.088 35.25 ;
      RECT -20 -20 23.134 35.204 ;
      RECT -20 -20 23.18 35.158 ;
      RECT -20 -20 23.226 35.112 ;
      RECT -20 -20 23.272 35.066 ;
      RECT -20 -20 23.318 35.02 ;
      RECT -20 -20 23.364 34.974 ;
      RECT -20 -20 23.41 34.928 ;
      RECT -20 -20 23.456 34.882 ;
      RECT -20 -20 23.502 34.836 ;
      RECT -20 -20 23.548 34.79 ;
      RECT -20 -20 23.594 34.744 ;
      RECT -20 -20 23.64 34.698 ;
      RECT -20 -20 23.686 34.652 ;
      RECT -20 -20 23.732 34.606 ;
      RECT -20 -20 23.778 34.56 ;
      RECT -20 -20 23.824 34.514 ;
      RECT -20 -20 23.87 34.468 ;
      RECT -20 -20 23.916 34.422 ;
      RECT -20 -20 23.962 34.376 ;
      RECT -20 -20 24.008 34.33 ;
      RECT -20 -20 24.054 34.284 ;
      RECT -20 -20 24.1 34.238 ;
      RECT -20 -20 24.146 34.192 ;
      RECT -20 -20 24.192 34.146 ;
      RECT -20 -20 24.238 34.1 ;
      RECT -20 -20 24.284 34.054 ;
      RECT -20 -20 24.33 34.008 ;
      RECT -20 -20 24.376 33.962 ;
      RECT -20 -20 24.422 33.916 ;
      RECT -20 -20 24.468 33.87 ;
      RECT -20 -20 24.514 33.824 ;
      RECT -20 -20 24.56 33.778 ;
      RECT -20 -20 24.606 33.732 ;
      RECT -20 -20 24.652 33.686 ;
      RECT -20 -20 24.698 33.64 ;
      RECT -20 -20 24.744 33.594 ;
      RECT -20 -20 24.79 33.548 ;
      RECT -20 -20 24.836 33.502 ;
      RECT -20 -20 24.882 33.456 ;
      RECT -20 -20 24.928 33.41 ;
      RECT -20 -20 24.974 33.364 ;
      RECT -20 -20 25.02 33.318 ;
      RECT -20 -20 25.066 33.272 ;
      RECT -20 -20 25.112 33.226 ;
      RECT -20 -20 25.158 33.18 ;
      RECT -20 -20 25.204 33.134 ;
      RECT -20 -20 25.25 33.088 ;
      RECT -20 -20 25.296 33.042 ;
      RECT -20 -20 25.342 32.996 ;
      RECT -20 -20 25.388 32.95 ;
      RECT -20 -20 25.434 32.904 ;
      RECT -20 -20 25.48 32.858 ;
      RECT -20 -20 25.526 32.812 ;
      RECT -20 -20 25.572 32.766 ;
      RECT -20 -20 25.618 32.72 ;
      RECT -20 -20 25.664 32.674 ;
      RECT -20 -20 25.71 32.628 ;
      RECT -20 -20 25.756 32.582 ;
      RECT -20 -20 25.802 32.536 ;
      RECT -20 -20 25.848 32.49 ;
      RECT -20 -20 25.894 32.444 ;
      RECT -20 -20 25.94 32.398 ;
      RECT -20 -20 25.986 32.352 ;
      RECT -20 -20 26.032 32.306 ;
      RECT -20 -20 26.078 32.26 ;
      RECT -20 -20 26.124 32.214 ;
      RECT -20 -20 26.17 32.168 ;
      RECT -20 -20 26.216 32.122 ;
      RECT -20 -20 26.262 32.076 ;
      RECT -20 -20 26.308 32.03 ;
      RECT -20 -20 26.354 31.984 ;
      RECT -20 -20 26.4 31.938 ;
      RECT -20 -20 26.446 31.892 ;
      RECT -20 -20 26.492 31.846 ;
      RECT -20 -20 26.538 31.8 ;
      RECT -20 -20 26.584 31.754 ;
      RECT -20 -20 26.63 31.708 ;
      RECT -20 -20 26.676 31.662 ;
      RECT -20 -20 26.722 31.616 ;
      RECT -20 -20 26.768 31.57 ;
      RECT -20 -20 26.814 31.524 ;
      RECT -20 -20 26.86 31.478 ;
      RECT -20 -20 26.906 31.432 ;
      RECT -20 -20 26.952 31.386 ;
      RECT -20 -20 26.998 31.34 ;
      RECT -20 -20 27.044 31.294 ;
      RECT -20 -20 27.09 31.248 ;
      RECT -20 -20 27.136 31.202 ;
      RECT -20 -20 27.182 31.156 ;
      RECT -20 -20 27.228 31.11 ;
      RECT -20 -20 27.274 31.064 ;
      RECT -20 -20 27.32 31.018 ;
      RECT -20 -20 27.366 30.972 ;
      RECT -20 -20 27.412 30.926 ;
      RECT -20 -20 27.458 30.88 ;
      RECT -20 -20 27.504 30.834 ;
      RECT -20 -20 27.55 30.788 ;
      RECT -20 -20 27.596 30.742 ;
      RECT -20 -20 27.642 30.696 ;
      RECT -20 -20 27.688 30.65 ;
      RECT -20 -20 27.734 30.604 ;
      RECT -20 -20 27.78 30.558 ;
      RECT -20 -20 27.826 30.512 ;
      RECT -20 -20 27.872 30.466 ;
      RECT -20 -20 27.918 30.42 ;
      RECT -20 -20 27.964 30.374 ;
      RECT -20 -20 28.01 30.328 ;
      RECT -20 -20 28.056 30.282 ;
      RECT -20 -20 28.102 30.236 ;
      RECT -20 -20 28.148 30.19 ;
      RECT -20 -20 28.194 30.144 ;
      RECT -20 -20 28.24 30.098 ;
      RECT -20 -20 28.286 30.052 ;
      RECT -20 -20 28.332 30.006 ;
      RECT -20 -20 28.378 29.96 ;
      RECT -20 -20 28.424 29.914 ;
      RECT -20 -20 28.47 29.868 ;
      RECT -20 -20 28.516 29.822 ;
      RECT -20 -20 28.562 29.776 ;
      RECT -20 -20 28.608 29.73 ;
      RECT -20 -20 28.654 29.684 ;
      RECT -20 -20 28.7 29.638 ;
      RECT -20 -20 28.746 29.592 ;
      RECT -20 -20 28.792 29.546 ;
      RECT -20 -20 28.838 29.5 ;
      RECT -20 -20 28.884 29.454 ;
      RECT -20 -20 28.93 29.408 ;
      RECT -20 -20 28.976 29.362 ;
      RECT -20 -20 29.022 29.316 ;
      RECT -20 -20 29.068 29.27 ;
      RECT -20 -20 29.114 29.224 ;
      RECT -20 -20 29.16 29.178 ;
      RECT -20 -20 29.206 29.132 ;
      RECT -20 -20 29.252 29.086 ;
      RECT -20 -20 29.298 29.04 ;
      RECT -20 -20 29.344 28.994 ;
      RECT -20 -20 29.39 28.948 ;
      RECT -20 -20 29.436 28.902 ;
      RECT -20 -20 29.482 28.856 ;
      RECT -20 -20 29.528 28.81 ;
      RECT -20 -20 29.574 28.764 ;
      RECT -20 -20 29.62 28.718 ;
      RECT -20 -20 29.666 28.672 ;
      RECT -20 -20 29.712 28.626 ;
      RECT -20 -20 29.758 28.58 ;
      RECT -20 -20 29.804 28.534 ;
      RECT -20 -20 29.85 28.488 ;
      RECT -20 -20 29.896 28.442 ;
      RECT -20 -20 29.942 28.396 ;
      RECT -20 -20 29.988 28.35 ;
      RECT -20 -20 30.034 28.304 ;
      RECT -20 -20 30.08 28.258 ;
      RECT -20 -20 30.126 28.212 ;
      RECT -20 -20 30.172 28.166 ;
      RECT -20 -20 30.218 28.12 ;
      RECT -20 -20 30.264 28.074 ;
      RECT -20 -20 30.31 28.028 ;
      RECT -20 -20 30.356 27.982 ;
      RECT -20 -20 30.402 27.936 ;
      RECT -20 -20 30.448 27.89 ;
      RECT -20 -20 30.494 27.844 ;
      RECT -20 -20 30.54 27.798 ;
      RECT -20 -20 30.586 27.752 ;
      RECT -20 -20 30.632 27.706 ;
      RECT -20 -20 30.678 27.66 ;
      RECT -20 -20 30.724 27.614 ;
      RECT -20 -20 30.77 27.568 ;
      RECT -20 -20 30.816 27.522 ;
      RECT -20 -20 30.862 27.476 ;
      RECT -20 -20 30.908 27.43 ;
      RECT -20 -20 30.954 27.384 ;
      RECT -20 -20 31 27.338 ;
      RECT -20 -20 31.046 27.292 ;
      RECT -20 -20 31.092 27.246 ;
      RECT -20 -20 31.138 27.2 ;
      RECT -20 -20 31.184 27.154 ;
      RECT -20 -20 31.23 27.108 ;
      RECT -20 -20 31.276 27.062 ;
      RECT -20 -20 31.322 27.016 ;
      RECT -20 -20 31.368 26.97 ;
      RECT -20 -20 31.414 26.924 ;
      RECT -20 -20 31.46 26.878 ;
      RECT -20 -20 31.506 26.832 ;
      RECT -20 -20 31.552 26.786 ;
      RECT -20 -20 31.598 26.74 ;
      RECT -20 -20 31.644 26.694 ;
      RECT -20 -20 31.69 26.648 ;
      RECT -20 -20 31.736 26.602 ;
      RECT -20 -20 31.782 26.556 ;
      RECT -20 -20 31.828 26.51 ;
      RECT -20 -20 31.874 26.464 ;
      RECT -20 -20 31.92 26.418 ;
      RECT -20 -20 31.966 26.372 ;
      RECT -20 -20 32.012 26.326 ;
      RECT -20 -20 32.058 26.28 ;
      RECT -20 -20 32.104 26.234 ;
      RECT -20 -20 32.15 26.188 ;
      RECT -20 -20 32.196 26.142 ;
      RECT -20 -20 32.242 26.096 ;
      RECT -20 -20 32.288 26.05 ;
      RECT -20 -20 32.334 26.004 ;
      RECT -20 -20 32.38 25.958 ;
      RECT -20 -20 32.426 25.912 ;
      RECT -20 -20 32.472 25.866 ;
      RECT -20 -20 32.518 25.82 ;
      RECT -20 -20 32.564 25.774 ;
      RECT -20 -20 32.61 25.728 ;
      RECT -20 -20 32.656 25.682 ;
      RECT -20 -20 32.702 25.636 ;
      RECT -20 -20 32.748 25.59 ;
      RECT -20 -20 32.794 25.544 ;
      RECT -20 -20 32.84 25.498 ;
      RECT -20 -20 32.886 25.452 ;
      RECT -20 -20 32.932 25.406 ;
      RECT -20 -20 32.978 25.36 ;
      RECT -20 -20 33.024 25.314 ;
      RECT -20 -20 33.07 25.268 ;
      RECT -20 -20 33.116 25.222 ;
      RECT -20 -20 33.162 25.176 ;
      RECT -20 -20 33.208 25.13 ;
      RECT -20 -20 33.254 25.084 ;
      RECT -20 -20 33.3 25.038 ;
      RECT -20 -20 33.346 24.992 ;
      RECT -20 -20 33.392 24.946 ;
      RECT -20 -20 33.438 24.9 ;
      RECT -20 -20 33.484 24.854 ;
      RECT -20 -20 33.53 24.808 ;
      RECT -20 -20 33.576 24.762 ;
      RECT -20 -20 33.622 24.716 ;
      RECT -20 -20 33.668 24.67 ;
      RECT -20 -20 33.714 24.624 ;
      RECT -20 -20 33.76 24.578 ;
      RECT -20 -20 33.806 24.532 ;
      RECT -20 -20 33.852 24.486 ;
      RECT -20 -20 33.898 24.44 ;
      RECT -20 -20 33.944 24.394 ;
      RECT -20 -20 33.99 24.348 ;
      RECT -20 -20 34.036 24.302 ;
      RECT -20 -20 34.082 24.256 ;
      RECT -20 -20 34.128 24.21 ;
      RECT -20 -20 34.174 24.164 ;
      RECT -20 -20 34.22 24.118 ;
      RECT -20 -20 34.266 24.072 ;
      RECT -20 -20 34.312 24.026 ;
      RECT -20 -20 34.358 23.98 ;
      RECT -20 -20 34.404 23.934 ;
      RECT -20 -20 34.45 23.888 ;
      RECT -20 -20 34.496 23.842 ;
      RECT -20 -20 34.542 23.796 ;
      RECT -20 -20 34.588 23.75 ;
      RECT -20 -20 34.634 23.704 ;
      RECT -20 -20 34.68 23.658 ;
      RECT -20 -20 34.726 23.612 ;
      RECT -20 -20 34.772 23.566 ;
      RECT -20 -20 34.818 23.52 ;
      RECT -20 -20 34.864 23.474 ;
      RECT -20 -20 34.91 23.428 ;
      RECT -20 -20 34.956 23.382 ;
      RECT -20 -20 35.002 23.336 ;
      RECT -20 -20 35.048 23.29 ;
      RECT -20 -20 35.094 23.244 ;
      RECT -20 -20 35.14 23.198 ;
      RECT -20 -20 35.186 23.152 ;
      RECT -20 -20 35.232 23.106 ;
      RECT -20 -20 35.278 23.06 ;
      RECT -20 -20 35.324 23.014 ;
      RECT -20 -20 35.37 22.968 ;
      RECT -20 -20 35.416 22.922 ;
      RECT -20 -20 35.462 22.876 ;
      RECT -20 -20 35.508 22.83 ;
      RECT -20 -20 35.554 22.784 ;
      RECT -20 -20 35.6 22.738 ;
      RECT -20 -20 35.646 22.692 ;
      RECT -20 -20 35.692 22.646 ;
      RECT -20 -20 35.738 22.6 ;
      RECT -20 -20 35.784 22.554 ;
      RECT -20 -20 35.83 22.508 ;
      RECT -20 -20 35.876 22.462 ;
      RECT -20 -20 35.922 22.416 ;
      RECT -20 -20 35.968 22.37 ;
      RECT -20 -20 36.014 22.324 ;
      RECT -20 -20 36.06 22.278 ;
      RECT -20 -20 36.106 22.232 ;
      RECT -20 -20 36.152 22.186 ;
      RECT -20 -20 36.198 22.14 ;
      RECT -20 -20 36.244 22.094 ;
      RECT -20 -20 36.29 22.048 ;
      RECT -20 -20 36.336 22.002 ;
      RECT -20 -20 36.382 21.956 ;
      RECT -20 -20 36.428 21.91 ;
      RECT -20 -20 36.474 21.864 ;
      RECT -20 -20 36.52 21.818 ;
      RECT -20 -20 36.566 21.772 ;
      RECT -20 -20 36.612 21.726 ;
      RECT -20 -20 36.658 21.68 ;
      RECT -20 -20 36.704 21.634 ;
      RECT -20 -20 36.75 21.588 ;
      RECT -20 -20 36.796 21.542 ;
      RECT -20 -20 36.842 21.496 ;
      RECT -20 -20 36.888 21.45 ;
      RECT -20 -20 36.934 21.404 ;
      RECT -20 -20 36.98 21.358 ;
      RECT -20 -20 37.026 21.312 ;
      RECT -20 -20 37.072 21.266 ;
      RECT -20 -20 37.118 21.22 ;
      RECT -20 -20 37.164 21.174 ;
      RECT -20 -20 37.21 21.128 ;
      RECT -20 -20 37.256 21.082 ;
      RECT -20 -20 37.302 21.036 ;
      RECT -20 -20 37.348 20.99 ;
      RECT -20 -20 37.394 20.944 ;
      RECT -20 -20 37.44 20.898 ;
      RECT -20 -20 37.486 20.852 ;
      RECT -20 -20 37.532 20.806 ;
      RECT -20 -20 37.578 20.76 ;
      RECT -20 -20 37.624 20.714 ;
      RECT -20 -20 37.67 20.668 ;
      RECT -20 -20 37.716 20.622 ;
      RECT -20 -20 37.762 20.576 ;
      RECT -20 -20 37.808 20.53 ;
      RECT -20 -20 37.854 20.484 ;
      RECT -20 -20 37.9 20.438 ;
      RECT -20 -20 37.946 20.392 ;
      RECT -20 -20 37.992 20.346 ;
      RECT -20 -20 38.038 20.3 ;
      RECT -20 -20 38.084 20.254 ;
      RECT -20 -20 38.13 20.208 ;
      RECT -20 -20 38.176 20.162 ;
      RECT -20 -20 38.222 20.116 ;
      RECT -20 -20 38.268 20.07 ;
      RECT -20 -20 38.314 20.024 ;
      RECT -20 -20 38.36 19.978 ;
      RECT -20 -20 38.406 19.932 ;
      RECT -20 -20 38.452 19.886 ;
      RECT -20 -20 38.498 19.84 ;
      RECT -20 -20 38.544 19.794 ;
      RECT -20 -20 38.59 19.748 ;
      RECT -20 -20 38.636 19.702 ;
      RECT -20 -20 38.682 19.656 ;
      RECT -20 -20 38.728 19.61 ;
      RECT -20 -20 38.774 19.564 ;
      RECT -20 -20 38.82 19.518 ;
      RECT -20 -20 38.866 19.472 ;
      RECT -20 -20 38.912 19.426 ;
      RECT -20 -20 38.958 19.38 ;
      RECT -20 -20 39.004 19.334 ;
      RECT -20 -20 39.05 19.288 ;
      RECT -20 -20 39.096 19.242 ;
      RECT -20 -20 39.142 19.196 ;
      RECT -20 -20 39.188 19.15 ;
      RECT -20 -20 39.234 19.104 ;
      RECT -20 -20 39.28 19.058 ;
      RECT -20 -20 39.326 19.012 ;
      RECT -20 -20 39.372 18.966 ;
      RECT -20 -20 39.418 18.92 ;
      RECT -20 -20 39.464 18.874 ;
      RECT -20 -20 39.51 18.828 ;
      RECT -20 -20 39.556 18.782 ;
      RECT -20 -20 39.602 18.736 ;
      RECT -20 -20 39.648 18.69 ;
      RECT -20 -20 39.694 18.644 ;
      RECT -20 -20 39.74 18.598 ;
      RECT -20 -20 39.786 18.552 ;
      RECT -20 -20 39.832 18.506 ;
      RECT -20 -20 39.878 18.46 ;
      RECT -20 -20 39.924 18.414 ;
      RECT -20 -20 39.97 18.368 ;
      RECT -20 -20 40.016 18.322 ;
      RECT -20 -20 40.062 18.276 ;
      RECT -20 -20 40.108 18.23 ;
      RECT -20 -20 40.154 18.184 ;
      RECT -20 -20 40.2 18.138 ;
      RECT -20 -20 40.246 18.092 ;
      RECT -20 -20 40.292 18.046 ;
      RECT -20 -20 40.338 18 ;
      RECT -20 -20 40.384 17.954 ;
      RECT -20 -20 40.43 17.908 ;
      RECT -20 -20 40.476 17.862 ;
      RECT -20 -20 40.522 17.816 ;
      RECT -20 -20 40.568 17.77 ;
      RECT -20 -20 40.614 17.724 ;
      RECT -20 -20 40.66 17.678 ;
      RECT -20 -20 40.706 17.632 ;
      RECT -20 -20 40.752 17.586 ;
      RECT -20 -20 40.798 17.54 ;
      RECT -20 -20 40.844 17.494 ;
      RECT -20 -20 40.89 17.448 ;
      RECT -20 -20 40.936 17.402 ;
      RECT -20 -20 40.982 17.356 ;
      RECT -20 -20 41.028 17.31 ;
      RECT -20 -20 41.074 17.264 ;
      RECT -20 -20 41.12 17.218 ;
      RECT -20 -20 41.166 17.172 ;
      RECT -20 -20 41.212 17.126 ;
      RECT -20 -20 41.258 17.08 ;
      RECT -20 -20 41.304 17.034 ;
      RECT -20 -20 41.35 16.988 ;
      RECT -20 -20 41.396 16.942 ;
      RECT -20 -20 41.442 16.896 ;
      RECT -20 -20 41.488 16.85 ;
      RECT -20 -20 41.534 16.804 ;
      RECT -20 -20 41.58 16.758 ;
      RECT -20 -20 41.626 16.712 ;
      RECT -20 -20 41.672 16.666 ;
      RECT -20 -20 41.718 16.62 ;
      RECT -20 -20 41.764 16.574 ;
      RECT -20 -20 41.81 16.528 ;
      RECT -20 -20 41.856 16.482 ;
      RECT -20 -20 41.902 16.436 ;
      RECT -20 -20 41.948 16.39 ;
      RECT -20 -20 41.994 16.344 ;
      RECT -20 -20 42.04 16.298 ;
      RECT -20 -20 42.086 16.252 ;
      RECT -20 -20 42.132 16.206 ;
      RECT -20 -20 42.178 16.16 ;
      RECT -20 -20 42.224 16.114 ;
      RECT -20 -20 42.27 16.068 ;
      RECT -20 -20 42.316 16.022 ;
      RECT -20 -20 42.362 15.976 ;
      RECT -20 -20 42.408 15.93 ;
      RECT -20 -20 42.454 15.884 ;
      RECT -20 -20 42.5 15.838 ;
      RECT -20 -20 42.546 15.792 ;
      RECT -20 -20 42.592 15.746 ;
      RECT -20 -20 42.638 15.7 ;
      RECT -20 -20 42.684 15.654 ;
      RECT -20 -20 42.73 15.608 ;
      RECT -20 -20 42.776 15.562 ;
      RECT -20 -20 42.822 15.516 ;
      RECT -20 -20 42.868 15.47 ;
      RECT -20 -20 42.914 15.424 ;
      RECT -20 -20 42.96 15.378 ;
      RECT -20 -20 43.006 15.332 ;
      RECT -20 -20 43.052 15.286 ;
      RECT -20 -20 43.098 15.24 ;
      RECT -20 -20 43.144 15.194 ;
      RECT -20 -20 43.19 15.148 ;
      RECT -20 -20 43.236 15.102 ;
      RECT -20 -20 43.282 15.056 ;
      RECT -20 -20 43.328 15.01 ;
      RECT -20 -20 43.374 14.964 ;
      RECT -20 -20 43.42 14.918 ;
      RECT -20 -20 43.466 14.872 ;
      RECT -20 -20 43.512 14.826 ;
      RECT -20 -20 43.558 14.78 ;
      RECT -20 -20 43.604 14.734 ;
      RECT -20 -20 43.65 14.688 ;
      RECT -20 -20 43.696 14.642 ;
      RECT -20 -20 43.742 14.596 ;
      RECT -20 -20 43.788 14.55 ;
      RECT -20 -20 43.834 14.504 ;
      RECT -20 -20 43.88 14.458 ;
      RECT -20 -20 43.926 14.412 ;
      RECT -20 -20 43.972 14.366 ;
      RECT -20 -20 44.018 14.32 ;
      RECT -20 -20 44.064 14.274 ;
      RECT -20 -20 44.11 14.228 ;
      RECT -20 -20 44.156 14.182 ;
      RECT -20 -20 44.202 14.136 ;
      RECT -20 -20 44.248 14.09 ;
      RECT -20 -20 44.294 14.044 ;
      RECT -20 -20 44.34 13.998 ;
      RECT -20 -20 44.386 13.952 ;
      RECT -20 -20 44.432 13.906 ;
      RECT -20 -20 44.478 13.86 ;
      RECT -20 -20 44.524 13.814 ;
      RECT -20 -20 44.57 13.768 ;
      RECT -20 -20 44.616 13.722 ;
      RECT -20 -20 44.662 13.676 ;
      RECT -20 -20 44.708 13.63 ;
      RECT -20 -20 44.754 13.584 ;
      RECT -20 -20 44.8 13.538 ;
      RECT -20 -20 44.846 13.492 ;
      RECT -20 -20 44.892 13.446 ;
      RECT -20 -20 44.938 13.4 ;
      RECT -20 -20 44.984 13.354 ;
      RECT -20 -20 45.03 13.308 ;
      RECT -20 -20 45.076 13.262 ;
      RECT -20 -20 45.122 13.216 ;
      RECT -20 -20 45.168 13.17 ;
      RECT -20 -20 45.214 13.124 ;
      RECT -20 -20 45.26 13.078 ;
      RECT -20 -20 45.306 13.032 ;
      RECT -20 -20 45.352 12.986 ;
      RECT -20 -20 45.398 12.94 ;
      RECT -20 -20 45.444 12.894 ;
      RECT -20 -20 45.49 12.848 ;
      RECT -20 -20 45.536 12.802 ;
      RECT -20 -20 45.582 12.756 ;
      RECT -20 -20 45.628 12.71 ;
      RECT -20 -20 45.674 12.664 ;
      RECT -20 -20 45.72 12.618 ;
      RECT -20 -20 45.766 12.572 ;
      RECT -20 -20 45.812 12.526 ;
      RECT -20 -20 45.858 12.48 ;
      RECT -20 -20 45.904 12.434 ;
      RECT -20 -20 45.95 12.388 ;
      RECT -20 -20 45.996 12.342 ;
      RECT -20 -20 46.042 12.296 ;
      RECT -20 -20 46.088 12.25 ;
      RECT -20 -20 46.134 12.204 ;
      RECT -20 -20 46.18 12.158 ;
      RECT -20 -20 46.226 12.112 ;
      RECT -20 -20 46.272 12.066 ;
      RECT -20 -20 46.318 12.02 ;
      RECT -20 -20 46.364 11.974 ;
      RECT -20 -20 46.41 11.928 ;
      RECT -20 -20 46.456 11.882 ;
      RECT -20 -20 46.502 11.836 ;
      RECT -20 -20 46.548 11.79 ;
      RECT -20 -20 46.594 11.744 ;
      RECT -20 -20 46.64 11.698 ;
      RECT -20 -20 46.686 11.652 ;
      RECT -20 -20 46.732 11.606 ;
      RECT -20 -20 46.778 11.56 ;
      RECT -20 -20 46.824 11.514 ;
      RECT -20 -20 46.87 11.468 ;
      RECT -20 -20 46.916 11.422 ;
      RECT -20 -20 46.962 11.376 ;
      RECT -20 -20 47.008 11.33 ;
      RECT -20 -20 47.054 11.284 ;
      RECT -20 -20 47.1 11.238 ;
      RECT -20 -20 47.146 11.192 ;
      RECT -20 -20 47.192 11.146 ;
      RECT -20 -20 47.238 11.1 ;
      RECT -20 -20 47.284 11.054 ;
      RECT -20 -20 47.33 11.008 ;
      RECT -20 -20 47.376 10.962 ;
      RECT -20 -20 47.422 10.916 ;
      RECT -20 -20 47.468 10.87 ;
      RECT -20 -20 47.514 10.824 ;
      RECT -20 -20 47.56 10.778 ;
      RECT -20 -20 47.606 10.732 ;
      RECT -20 -20 47.652 10.686 ;
      RECT -20 -20 47.698 10.64 ;
      RECT -20 -20 47.744 10.594 ;
      RECT -20 -20 47.79 10.548 ;
      RECT -20 -20 47.836 10.502 ;
      RECT -20 -20 47.882 10.456 ;
      RECT -20 -20 47.928 10.41 ;
      RECT -20 -20 47.974 10.364 ;
      RECT -20 -20 48.02 10.318 ;
      RECT -20 -20 48.066 10.272 ;
      RECT -20 -20 48.112 10.226 ;
      RECT -20 -20 48.158 10.18 ;
      RECT -20 -20 48.204 10.134 ;
      RECT -20 -20 48.25 10.088 ;
      RECT -20 -20 48.296 10.042 ;
      RECT -20 -20 48.342 9.996 ;
      RECT -20 -20 48.388 9.95 ;
      RECT -20 -20 48.434 9.904 ;
      RECT -20 -20 48.48 9.858 ;
      RECT -20 -20 48.526 9.812 ;
      RECT -20 -20 48.572 9.766 ;
      RECT -20 -20 48.618 9.72 ;
      RECT -20 -20 48.664 9.674 ;
      RECT -20 -20 48.71 9.628 ;
      RECT -20 -20 48.756 9.582 ;
      RECT -20 -20 48.802 9.536 ;
      RECT -20 -20 48.848 9.49 ;
      RECT -20 -20 48.894 9.444 ;
      RECT -20 -20 48.94 9.398 ;
      RECT -20 -20 48.986 9.352 ;
      RECT -20 -20 49.032 9.306 ;
      RECT -20 -20 49.078 9.26 ;
      RECT -20 -20 49.124 9.214 ;
      RECT -20 -20 49.17 9.168 ;
      RECT -20 -20 49.216 9.122 ;
      RECT -20 -20 49.262 9.076 ;
      RECT -20 -20 49.308 9.03 ;
      RECT -20 -20 49.354 8.984 ;
      RECT -20 -20 49.4 8.938 ;
      RECT -20 -20 49.446 8.892 ;
      RECT -20 -20 49.492 8.846 ;
      RECT -20 -20 49.538 8.8 ;
      RECT -20 -20 49.584 8.754 ;
      RECT -20 -20 49.63 8.708 ;
      RECT -20 -20 49.676 8.662 ;
      RECT -20 -20 49.722 8.616 ;
      RECT -20 -20 49.768 8.57 ;
      RECT -20 -20 49.814 8.524 ;
      RECT -20 -20 49.86 8.478 ;
      RECT -20 -20 49.906 8.432 ;
      RECT -20 -20 49.952 8.386 ;
      RECT -20 -20 49.998 8.34 ;
      RECT -20 -20 50.044 8.294 ;
      RECT -20 -20 50.09 8.248 ;
      RECT -20 -20 50.136 8.202 ;
      RECT -20 -20 50.182 8.156 ;
      RECT -20 -20 50.228 8.11 ;
      RECT -20 -20 50.274 8.064 ;
      RECT -20 -20 50.32 8.018 ;
      RECT -20 -20 50.366 7.972 ;
      RECT -20 -20 50.412 7.926 ;
      RECT -20 -20 50.458 7.88 ;
      RECT -20 -20 50.504 7.834 ;
      RECT -20 -20 50.55 7.788 ;
      RECT -20 -20 50.596 7.742 ;
      RECT -20 -20 50.642 7.696 ;
      RECT -20 -20 50.688 7.65 ;
      RECT -20 -20 50.734 7.604 ;
      RECT -20 -20 50.78 7.558 ;
      RECT -20 -20 50.826 7.512 ;
      RECT -20 -20 50.872 7.466 ;
      RECT -20 -20 50.918 7.42 ;
      RECT -20 -20 50.964 7.374 ;
      RECT -20 -20 51.01 7.328 ;
      RECT -20 -20 51.056 7.282 ;
      RECT -20 -20 51.102 7.236 ;
      RECT -20 -20 51.148 7.19 ;
      RECT -20 -20 51.194 7.144 ;
      RECT -20 -20 51.24 7.098 ;
      RECT -20 -20 51.286 7.052 ;
      RECT -20 -20 51.332 7.006 ;
      RECT -20 -20 51.378 6.96 ;
      RECT -20 -20 51.424 6.914 ;
      RECT -20 -20 51.47 6.868 ;
      RECT -20 -20 51.516 6.822 ;
      RECT -20 -20 51.562 6.776 ;
      RECT -20 -20 51.608 6.73 ;
      RECT -20 -20 51.654 6.684 ;
      RECT -20 -20 51.7 6.638 ;
      RECT -20 -20 51.746 6.592 ;
      RECT -20 -20 51.792 6.546 ;
      RECT -20 -20 51.838 6.5 ;
      RECT -20 -20 51.884 6.454 ;
      RECT -20 -20 51.93 6.408 ;
      RECT -20 -20 51.976 6.362 ;
      RECT -20 -20 52.022 6.316 ;
      RECT -20 -20 52.068 6.27 ;
      RECT -20 -20 52.114 6.224 ;
      RECT -20 -20 52.16 6.178 ;
      RECT -20 -20 52.206 6.132 ;
      RECT -20 -20 52.252 6.086 ;
      RECT -20 -20 52.298 6.04 ;
      RECT -20 -20 52.344 5.994 ;
      RECT -20 -20 52.39 5.948 ;
      RECT -20 -20 52.436 5.902 ;
      RECT -20 -20 52.482 5.856 ;
      RECT -20 -20 52.528 5.81 ;
      RECT -20 -20 52.574 5.764 ;
      RECT -20 -20 52.62 5.718 ;
      RECT -20 -20 52.666 5.672 ;
      RECT -20 -20 52.712 5.626 ;
      RECT -20 -20 52.758 5.58 ;
      RECT -20 -20 52.804 5.534 ;
      RECT -20 -20 52.85 5.488 ;
      RECT -20 -20 52.896 5.442 ;
      RECT -20 -20 52.942 5.396 ;
      RECT -20 -20 52.988 5.35 ;
      RECT -20 -20 53.034 5.304 ;
      RECT -20 -20 53.08 5.258 ;
      RECT -20 -20 53.126 5.212 ;
      RECT -20 -20 53.172 5.166 ;
      RECT -20 -20 53.218 5.12 ;
      RECT -20 -20 53.264 5.074 ;
      RECT -20 -20 53.31 5.028 ;
      RECT -20 -20 53.356 4.982 ;
      RECT -20 -20 53.402 4.936 ;
      RECT -20 -20 53.448 4.89 ;
      RECT -20 -20 53.494 4.844 ;
      RECT -20 -20 53.54 4.798 ;
      RECT -20 -20 53.586 4.752 ;
      RECT -20 -20 53.632 4.706 ;
      RECT -20 -20 53.678 4.66 ;
      RECT -20 -20 53.724 4.614 ;
      RECT -20 -20 53.77 4.568 ;
      RECT -20 -20 53.816 4.522 ;
      RECT -20 -20 53.862 4.476 ;
      RECT -20 -20 53.908 4.43 ;
      RECT -20 -20 53.954 4.384 ;
      RECT -20 -20 54 4.338 ;
      RECT -20 -20 54.046 4.292 ;
      RECT -20 -20 54.092 4.246 ;
      RECT -20 -20 54.138 4.2 ;
      RECT -20 -20 54.184 4.154 ;
      RECT -20 -20 54.23 4.108 ;
      RECT -20 -20 54.276 4.062 ;
      RECT -20 -20 54.322 4.016 ;
      RECT -20 -20 54.368 3.97 ;
      RECT -20 -20 54.414 3.924 ;
      RECT -20 -20 54.46 3.878 ;
      RECT -20 -20 54.506 3.832 ;
      RECT -20 -20 54.552 3.786 ;
      RECT -20 -20 54.598 3.74 ;
      RECT -20 -20 54.644 3.694 ;
      RECT -20 -20 54.69 3.648 ;
      RECT -20 -20 54.736 3.602 ;
      RECT -20 -20 54.782 3.556 ;
      RECT -20 -20 54.828 3.51 ;
      RECT -20 -20 54.874 3.464 ;
      RECT -20 -20 54.92 3.418 ;
      RECT -20 -20 54.966 3.372 ;
      RECT -20 -20 55.012 3.326 ;
      RECT -20 -20 55.058 3.28 ;
      RECT -20 -20 55.104 3.234 ;
      RECT -20 -20 55.15 3.188 ;
      RECT -20 -20 55.196 3.142 ;
      RECT -20 -20 55.242 3.096 ;
      RECT -20 -20 55.288 3.05 ;
      RECT -20 -20 55.334 3.004 ;
      RECT -20 -20 55.38 2.958 ;
      RECT -20 -20 55.415 2.917 ;
      RECT -20 -20 110 2.9 ;
      RECT 64.1 85.817 67.9 110 ;
      RECT 64.1 85.817 67.946 87.742 ;
      RECT 64.1 85.817 67.992 87.696 ;
      RECT 64.1 85.817 68.038 87.65 ;
      RECT 64.1 85.817 68.084 87.604 ;
      RECT 64.1 85.817 68.13 87.558 ;
      RECT 64.1 85.817 68.176 87.512 ;
      RECT 64.1 85.817 68.222 87.466 ;
      RECT 64.1 85.817 68.268 87.42 ;
      RECT 64.1 85.817 68.314 87.374 ;
      RECT 64.1 85.817 68.36 87.328 ;
      RECT 64.1 85.817 68.406 87.282 ;
      RECT 64.1 85.817 68.452 87.236 ;
      RECT 64.1 85.817 68.498 87.19 ;
      RECT 64.1 85.817 68.544 87.144 ;
      RECT 64.1 85.817 68.59 87.098 ;
      RECT 64.1 85.817 68.636 87.052 ;
      RECT 64.1 85.817 68.682 87.006 ;
      RECT 64.1 85.817 68.728 86.96 ;
      RECT 64.1 85.817 68.774 86.914 ;
      RECT 64.1 85.817 68.82 86.868 ;
      RECT 64.1 85.817 68.866 86.822 ;
      RECT 64.1 85.817 68.912 86.776 ;
      RECT 64.1 85.817 68.958 86.73 ;
      RECT 64.1 85.817 69.004 86.684 ;
      RECT 64.1 85.817 69.05 86.638 ;
      RECT 64.1 85.817 69.096 86.592 ;
      RECT 64.1 85.817 69.142 86.546 ;
      RECT 64.1 85.817 69.188 86.5 ;
      RECT 64.1 85.817 69.234 86.454 ;
      RECT 64.1 85.817 69.28 86.408 ;
      RECT 64.1 85.817 69.326 86.362 ;
      RECT 64.1 85.817 69.372 86.316 ;
      RECT 64.1 85.817 69.418 86.27 ;
      RECT 64.1 85.817 69.464 86.224 ;
      RECT 64.1 85.817 69.51 86.178 ;
      RECT 64.1 85.817 69.556 86.132 ;
      RECT 64.1 85.817 69.602 86.086 ;
      RECT 64.1 85.817 69.648 86.04 ;
      RECT 64.1 85.817 69.694 85.994 ;
      RECT 64.1 85.817 69.74 85.948 ;
      RECT 64.1 85.817 69.786 85.902 ;
      RECT 64.146 85.771 69.832 85.856 ;
      RECT 64.192 85.725 69.878 85.81 ;
      RECT 64.238 85.679 69.924 85.764 ;
      RECT 64.284 85.633 69.97 85.718 ;
      RECT 64.33 85.587 70.016 85.672 ;
      RECT 64.376 85.541 70.062 85.626 ;
      RECT 64.422 85.495 70.108 85.58 ;
      RECT 64.468 85.449 70.154 85.534 ;
      RECT 64.514 85.403 70.2 85.488 ;
      RECT 64.56 85.357 70.246 85.442 ;
      RECT 64.606 85.311 70.292 85.396 ;
      RECT 64.652 85.265 70.338 85.35 ;
      RECT 64.698 85.219 70.384 85.304 ;
      RECT 64.744 85.173 70.43 85.258 ;
      RECT 64.79 85.127 70.476 85.212 ;
      RECT 64.836 85.081 70.522 85.166 ;
      RECT 64.882 85.035 70.568 85.12 ;
      RECT 64.928 84.989 70.614 85.074 ;
      RECT 64.974 84.943 70.66 85.028 ;
      RECT 65.02 84.897 70.706 84.982 ;
      RECT 65.066 84.851 70.752 84.936 ;
      RECT 65.112 84.805 70.798 84.89 ;
      RECT 65.158 84.759 70.844 84.844 ;
      RECT 65.204 84.713 70.89 84.798 ;
      RECT 65.25 84.667 70.936 84.752 ;
      RECT 65.296 84.621 70.982 84.706 ;
      RECT 65.342 84.575 71.028 84.66 ;
      RECT 65.388 84.529 71.074 84.614 ;
      RECT 65.434 84.483 71.12 84.568 ;
      RECT 65.48 84.437 71.166 84.522 ;
      RECT 65.526 84.391 71.212 84.476 ;
      RECT 65.572 84.345 71.258 84.43 ;
      RECT 65.618 84.299 71.304 84.384 ;
      RECT 65.664 84.253 71.35 84.338 ;
      RECT 65.71 84.207 71.396 84.292 ;
      RECT 65.756 84.161 71.442 84.246 ;
      RECT 65.802 84.115 71.488 84.2 ;
      RECT 65.848 84.069 71.534 84.154 ;
      RECT 65.894 84.023 71.58 84.108 ;
      RECT 65.94 83.977 71.626 84.062 ;
      RECT 65.986 83.931 71.672 84.016 ;
      RECT 66.032 83.885 71.718 83.97 ;
      RECT 66.078 83.839 71.764 83.924 ;
      RECT 66.124 83.793 71.81 83.878 ;
      RECT 66.17 83.747 71.856 83.832 ;
      RECT 66.216 83.701 71.902 83.786 ;
      RECT 66.262 83.655 71.948 83.74 ;
      RECT 66.308 83.609 71.994 83.694 ;
      RECT 66.354 83.563 72.04 83.648 ;
      RECT 66.4 83.517 72.086 83.602 ;
      RECT 66.446 83.471 72.132 83.556 ;
      RECT 66.492 83.425 72.178 83.51 ;
      RECT 66.538 83.379 72.224 83.464 ;
      RECT 66.584 83.333 72.27 83.418 ;
      RECT 66.63 83.287 72.316 83.372 ;
      RECT 66.676 83.241 72.362 83.326 ;
      RECT 66.722 83.195 72.408 83.28 ;
      RECT 66.768 83.149 72.454 83.234 ;
      RECT 66.814 83.103 72.5 83.188 ;
      RECT 66.86 83.057 72.546 83.142 ;
      RECT 66.906 83.011 72.592 83.096 ;
      RECT 66.952 82.965 72.638 83.05 ;
      RECT 66.998 82.919 72.684 83.004 ;
      RECT 67.044 82.873 72.73 82.958 ;
      RECT 67.09 82.827 72.776 82.912 ;
      RECT 67.136 82.781 72.822 82.866 ;
      RECT 67.182 82.735 72.868 82.82 ;
      RECT 67.228 82.689 72.914 82.774 ;
      RECT 67.274 82.643 72.96 82.728 ;
      RECT 67.32 82.597 73.006 82.682 ;
      RECT 67.366 82.551 73.052 82.636 ;
      RECT 67.412 82.505 73.098 82.59 ;
      RECT 67.458 82.459 73.144 82.544 ;
      RECT 67.504 82.413 73.19 82.498 ;
      RECT 67.55 82.367 73.236 82.452 ;
      RECT 67.596 82.321 73.282 82.406 ;
      RECT 67.642 82.275 73.328 82.36 ;
      RECT 67.688 82.229 73.374 82.314 ;
      RECT 67.734 82.183 73.42 82.268 ;
      RECT 67.78 82.137 73.466 82.222 ;
      RECT 67.826 82.091 73.512 82.176 ;
      RECT 67.872 82.045 73.558 82.13 ;
      RECT 67.918 81.999 73.604 82.084 ;
      RECT 67.964 81.953 73.65 82.038 ;
      RECT 68.01 81.907 73.696 81.992 ;
      RECT 68.056 81.861 73.742 81.946 ;
      RECT 68.102 81.815 73.788 81.9 ;
      RECT 68.148 81.769 73.834 81.854 ;
      RECT 68.194 81.723 73.88 81.808 ;
      RECT 68.24 81.677 73.926 81.762 ;
      RECT 68.286 81.631 73.972 81.716 ;
      RECT 68.332 81.585 74.018 81.67 ;
      RECT 68.378 81.539 74.064 81.624 ;
      RECT 68.424 81.493 74.11 81.578 ;
      RECT 68.47 81.447 74.156 81.532 ;
      RECT 68.516 81.401 74.202 81.486 ;
      RECT 68.562 81.355 74.248 81.44 ;
      RECT 68.608 81.309 74.294 81.394 ;
      RECT 68.654 81.263 74.34 81.348 ;
      RECT 68.7 81.217 74.386 81.302 ;
      RECT 68.746 81.171 74.432 81.256 ;
      RECT 68.792 81.125 74.478 81.21 ;
      RECT 68.838 81.079 74.524 81.164 ;
      RECT 68.884 81.033 74.57 81.118 ;
      RECT 68.93 80.987 74.616 81.072 ;
      RECT 68.976 80.941 74.662 81.026 ;
      RECT 69.022 80.895 74.708 80.98 ;
      RECT 69.068 80.849 74.754 80.934 ;
      RECT 69.114 80.803 74.8 80.888 ;
      RECT 69.16 80.757 74.846 80.842 ;
      RECT 69.206 80.711 74.892 80.796 ;
      RECT 69.252 80.665 74.938 80.75 ;
      RECT 69.298 80.619 74.984 80.704 ;
      RECT 69.344 80.573 75.03 80.658 ;
      RECT 69.39 80.527 75.076 80.612 ;
      RECT 69.436 80.481 75.122 80.566 ;
      RECT 69.482 80.435 75.168 80.52 ;
      RECT 69.528 80.389 75.214 80.474 ;
      RECT 69.574 80.343 75.26 80.428 ;
      RECT 69.62 80.297 75.306 80.382 ;
      RECT 69.666 80.251 75.352 80.336 ;
      RECT 69.712 80.205 75.398 80.29 ;
      RECT 69.758 80.159 75.444 80.244 ;
      RECT 69.804 80.113 75.49 80.198 ;
      RECT 69.85 80.067 75.536 80.152 ;
      RECT 69.896 80.021 75.582 80.106 ;
      RECT 69.942 79.975 75.628 80.06 ;
      RECT 69.988 79.929 75.674 80.014 ;
      RECT 70.034 79.883 75.72 79.968 ;
      RECT 70.08 79.837 75.766 79.922 ;
      RECT 70.126 79.791 75.812 79.876 ;
      RECT 70.172 79.745 75.858 79.83 ;
      RECT 70.218 79.699 75.904 79.784 ;
      RECT 70.264 79.653 75.95 79.738 ;
      RECT 70.31 79.607 75.996 79.692 ;
      RECT 70.356 79.561 76.042 79.646 ;
      RECT 70.402 79.515 76.088 79.6 ;
      RECT 70.448 79.469 76.134 79.554 ;
      RECT 70.494 79.423 76.18 79.508 ;
      RECT 70.54 79.377 76.226 79.462 ;
      RECT 70.586 79.331 76.272 79.416 ;
      RECT 70.632 79.285 76.318 79.37 ;
      RECT 70.678 79.239 76.364 79.324 ;
      RECT 70.678 79.239 76.4 79.283 ;
      RECT 70.724 79.193 76.446 79.242 ;
      RECT 76.382 73.535 76.446 79.242 ;
      RECT 70.77 79.147 76.492 79.196 ;
      RECT 76.428 73.489 76.492 79.196 ;
      RECT 70.816 79.101 76.538 79.15 ;
      RECT 76.474 73.443 76.538 79.15 ;
      RECT 70.862 79.055 76.584 79.104 ;
      RECT 76.52 73.397 76.584 79.104 ;
      RECT 70.908 79.009 76.63 79.058 ;
      RECT 76.566 73.351 76.63 79.058 ;
      RECT 70.954 78.963 76.676 79.012 ;
      RECT 76.612 73.305 76.676 79.012 ;
      RECT 71 78.917 76.722 78.966 ;
      RECT 76.658 73.259 76.722 78.966 ;
      RECT 71.046 78.871 76.768 78.92 ;
      RECT 76.704 73.213 76.768 78.92 ;
      RECT 71.092 78.825 76.814 78.874 ;
      RECT 76.75 73.167 76.814 78.874 ;
      RECT 71.138 78.779 76.86 78.828 ;
      RECT 76.796 73.121 76.86 78.828 ;
      RECT 71.184 78.733 76.906 78.782 ;
      RECT 76.842 73.075 76.906 78.782 ;
      RECT 71.23 78.687 76.952 78.736 ;
      RECT 76.888 73.029 76.952 78.736 ;
      RECT 71.276 78.641 76.998 78.69 ;
      RECT 76.934 72.983 76.998 78.69 ;
      RECT 71.322 78.595 77.044 78.644 ;
      RECT 76.98 72.937 77.044 78.644 ;
      RECT 71.368 78.549 77.09 78.598 ;
      RECT 77.026 72.891 77.09 78.598 ;
      RECT 71.414 78.503 77.136 78.552 ;
      RECT 77.072 72.845 77.136 78.552 ;
      RECT 71.46 78.457 77.182 78.506 ;
      RECT 77.118 72.799 77.182 78.506 ;
      RECT 71.506 78.411 77.228 78.46 ;
      RECT 77.164 72.753 77.228 78.46 ;
      RECT 71.552 78.365 77.274 78.414 ;
      RECT 77.21 72.707 77.274 78.414 ;
      RECT 71.598 78.319 77.32 78.368 ;
      RECT 77.256 72.661 77.32 78.368 ;
      RECT 71.644 78.273 77.366 78.322 ;
      RECT 77.302 72.615 77.366 78.322 ;
      RECT 71.69 78.227 77.412 78.276 ;
      RECT 77.348 72.569 77.412 78.276 ;
      RECT 71.736 78.181 77.458 78.23 ;
      RECT 77.394 72.523 77.458 78.23 ;
      RECT 71.782 78.135 77.504 78.184 ;
      RECT 77.44 72.477 77.504 78.184 ;
      RECT 71.828 78.089 77.55 78.138 ;
      RECT 77.486 72.431 77.55 78.138 ;
      RECT 71.874 78.043 77.596 78.092 ;
      RECT 77.532 72.385 77.596 78.092 ;
      RECT 71.92 77.997 77.642 78.046 ;
      RECT 77.578 72.339 77.642 78.046 ;
      RECT 71.966 77.951 77.688 78 ;
      RECT 77.624 72.293 77.688 78 ;
      RECT 72.012 77.905 77.734 77.954 ;
      RECT 77.67 72.247 77.734 77.954 ;
      RECT 72.058 77.859 77.78 77.908 ;
      RECT 77.716 72.201 77.78 77.908 ;
      RECT 72.104 77.813 77.826 77.862 ;
      RECT 77.762 72.155 77.826 77.862 ;
      RECT 72.15 77.767 77.872 77.816 ;
      RECT 77.808 72.109 77.872 77.816 ;
      RECT 72.196 77.721 77.918 77.77 ;
      RECT 77.854 72.063 77.918 77.77 ;
      RECT 72.242 77.675 77.964 77.724 ;
      RECT 77.9 72.017 77.964 77.724 ;
      RECT 72.288 77.629 78.01 77.678 ;
      RECT 77.946 71.971 78.01 77.678 ;
      RECT 72.334 77.583 78.056 77.632 ;
      RECT 77.992 71.925 78.056 77.632 ;
      RECT 72.38 77.537 78.102 77.586 ;
      RECT 78.038 71.879 78.102 77.586 ;
      RECT 72.426 77.491 78.148 77.54 ;
      RECT 78.084 71.833 78.148 77.54 ;
      RECT 72.472 77.445 78.194 77.494 ;
      RECT 78.13 71.787 78.194 77.494 ;
      RECT 72.518 77.399 78.24 77.448 ;
      RECT 78.176 71.741 78.24 77.448 ;
      RECT 72.564 77.353 78.286 77.402 ;
      RECT 78.222 71.695 78.286 77.402 ;
      RECT 72.61 77.307 78.332 77.356 ;
      RECT 78.268 71.649 78.332 77.356 ;
      RECT 72.656 77.261 78.378 77.31 ;
      RECT 78.314 71.603 78.378 77.31 ;
      RECT 72.702 77.215 78.424 77.264 ;
      RECT 78.36 71.557 78.424 77.264 ;
      RECT 72.748 77.169 78.47 77.218 ;
      RECT 78.406 71.511 78.47 77.218 ;
      RECT 72.794 77.123 78.516 77.172 ;
      RECT 78.452 71.465 78.516 77.172 ;
      RECT 72.84 77.077 78.562 77.126 ;
      RECT 78.498 71.419 78.562 77.126 ;
      RECT 72.886 77.031 78.608 77.08 ;
      RECT 78.544 71.373 78.608 77.08 ;
      RECT 72.932 76.985 78.654 77.034 ;
      RECT 78.59 71.327 78.654 77.034 ;
      RECT 72.978 76.939 78.7 76.988 ;
      RECT 78.636 71.281 78.7 76.988 ;
      RECT 73.024 76.893 78.746 76.942 ;
      RECT 78.682 71.235 78.746 76.942 ;
      RECT 73.07 76.847 78.792 76.896 ;
      RECT 78.728 71.189 78.792 76.896 ;
      RECT 73.116 76.801 78.838 76.85 ;
      RECT 78.774 71.143 78.838 76.85 ;
      RECT 73.162 76.755 78.884 76.804 ;
      RECT 78.82 71.097 78.884 76.804 ;
      RECT 73.208 76.709 78.93 76.758 ;
      RECT 78.866 71.051 78.93 76.758 ;
      RECT 73.254 76.663 78.976 76.712 ;
      RECT 78.912 71.005 78.976 76.712 ;
      RECT 73.3 76.617 79.022 76.666 ;
      RECT 78.958 70.959 79.022 76.666 ;
      RECT 73.346 76.571 79.068 76.62 ;
      RECT 79.004 70.913 79.068 76.62 ;
      RECT 73.392 76.525 79.114 76.574 ;
      RECT 79.05 70.867 79.114 76.574 ;
      RECT 73.438 76.479 79.16 76.528 ;
      RECT 79.096 70.821 79.16 76.528 ;
      RECT 73.484 76.433 79.206 76.482 ;
      RECT 79.142 70.775 79.206 76.482 ;
      RECT 73.53 76.387 79.252 76.436 ;
      RECT 79.188 70.729 79.252 76.436 ;
      RECT 73.576 76.341 79.298 76.39 ;
      RECT 79.234 70.683 79.298 76.39 ;
      RECT 73.622 76.295 79.344 76.344 ;
      RECT 79.28 70.637 79.344 76.344 ;
      RECT 73.668 76.249 79.39 76.298 ;
      RECT 79.326 70.591 79.39 76.298 ;
      RECT 73.714 76.203 79.436 76.252 ;
      RECT 79.372 70.545 79.436 76.252 ;
      RECT 73.76 76.157 79.482 76.206 ;
      RECT 79.418 70.499 79.482 76.206 ;
      RECT 73.806 76.111 79.528 76.16 ;
      RECT 79.464 70.453 79.528 76.16 ;
      RECT 73.852 76.065 79.574 76.114 ;
      RECT 79.51 70.407 79.574 76.114 ;
      RECT 73.898 76.019 79.62 76.068 ;
      RECT 79.556 70.361 79.62 76.068 ;
      RECT 73.944 75.973 79.666 76.022 ;
      RECT 79.602 70.315 79.666 76.022 ;
      RECT 73.99 75.927 79.712 75.976 ;
      RECT 79.648 70.269 79.712 75.976 ;
      RECT 74.036 75.881 79.758 75.93 ;
      RECT 79.694 70.223 79.758 75.93 ;
      RECT 74.082 75.835 79.804 75.884 ;
      RECT 79.74 70.177 79.804 75.884 ;
      RECT 74.128 75.789 79.85 75.838 ;
      RECT 79.786 70.131 79.85 75.838 ;
      RECT 74.174 75.743 79.896 75.792 ;
      RECT 79.832 70.085 79.896 75.792 ;
      RECT 74.22 75.697 79.942 75.746 ;
      RECT 79.878 70.039 79.942 75.746 ;
      RECT 74.266 75.651 79.988 75.7 ;
      RECT 79.924 69.993 79.988 75.7 ;
      RECT 74.312 75.605 80.034 75.654 ;
      RECT 79.97 69.947 80.034 75.654 ;
      RECT 74.358 75.559 80.08 75.608 ;
      RECT 80.016 69.901 80.08 75.608 ;
      RECT 74.404 75.513 80.126 75.562 ;
      RECT 80.062 69.855 80.126 75.562 ;
      RECT 74.45 75.467 80.172 75.516 ;
      RECT 80.108 69.809 80.172 75.516 ;
      RECT 74.496 75.421 80.218 75.47 ;
      RECT 80.154 69.763 80.218 75.47 ;
      RECT 74.542 75.375 80.264 75.424 ;
      RECT 80.2 69.717 80.264 75.424 ;
      RECT 74.588 75.329 80.31 75.378 ;
      RECT 80.246 69.671 80.31 75.378 ;
      RECT 74.634 75.283 80.356 75.332 ;
      RECT 80.292 69.625 80.356 75.332 ;
      RECT 74.68 75.237 80.402 75.286 ;
      RECT 80.338 69.579 80.402 75.286 ;
      RECT 74.726 75.191 80.448 75.24 ;
      RECT 80.384 69.533 80.448 75.24 ;
      RECT 74.772 75.145 80.494 75.194 ;
      RECT 80.43 69.487 80.494 75.194 ;
      RECT 74.818 75.099 80.54 75.148 ;
      RECT 80.476 69.441 80.54 75.148 ;
      RECT 74.864 75.053 80.586 75.102 ;
      RECT 80.522 69.395 80.586 75.102 ;
      RECT 74.91 75.007 80.632 75.056 ;
      RECT 80.568 69.349 80.632 75.056 ;
      RECT 74.956 74.961 80.678 75.01 ;
      RECT 80.614 69.303 80.678 75.01 ;
      RECT 75.002 74.915 80.724 74.964 ;
      RECT 80.66 69.257 80.724 74.964 ;
      RECT 75.048 74.869 80.77 74.918 ;
      RECT 80.706 69.211 80.77 74.918 ;
      RECT 75.094 74.823 80.816 74.872 ;
      RECT 80.752 69.165 80.816 74.872 ;
      RECT 75.14 74.777 80.862 74.826 ;
      RECT 80.798 69.119 80.862 74.826 ;
      RECT 75.186 74.731 80.908 74.78 ;
      RECT 80.844 69.073 80.908 74.78 ;
      RECT 75.232 74.685 80.954 74.734 ;
      RECT 80.89 69.027 80.954 74.734 ;
      RECT 75.278 74.639 81 74.688 ;
      RECT 80.936 68.981 81 74.688 ;
      RECT 75.324 74.593 81.046 74.642 ;
      RECT 80.982 68.935 81.046 74.642 ;
      RECT 75.37 74.547 81.092 74.596 ;
      RECT 81.028 68.889 81.092 74.596 ;
      RECT 75.416 74.501 81.138 74.55 ;
      RECT 81.074 68.843 81.138 74.55 ;
      RECT 75.462 74.455 81.184 74.504 ;
      RECT 81.12 68.797 81.184 74.504 ;
      RECT 75.508 74.409 81.23 74.458 ;
      RECT 81.166 68.751 81.23 74.458 ;
      RECT 75.554 74.363 81.276 74.412 ;
      RECT 81.212 68.705 81.276 74.412 ;
      RECT 75.6 74.317 81.322 74.366 ;
      RECT 81.258 68.659 81.322 74.366 ;
      RECT 75.646 74.271 81.368 74.32 ;
      RECT 81.304 68.613 81.368 74.32 ;
      RECT 75.692 74.225 81.414 74.274 ;
      RECT 81.35 68.567 81.414 74.274 ;
      RECT 75.738 74.179 81.46 74.228 ;
      RECT 81.396 68.521 81.46 74.228 ;
      RECT 75.784 74.133 81.506 74.182 ;
      RECT 81.442 68.475 81.506 74.182 ;
      RECT 75.83 74.087 81.552 74.136 ;
      RECT 81.488 68.429 81.552 74.136 ;
      RECT 75.876 74.041 81.598 74.09 ;
      RECT 81.534 68.383 81.598 74.09 ;
      RECT 75.922 73.995 81.644 74.044 ;
      RECT 81.58 68.337 81.644 74.044 ;
      RECT 75.968 73.949 81.69 73.998 ;
      RECT 81.626 68.291 81.69 73.998 ;
      RECT 76.014 73.903 81.736 73.952 ;
      RECT 81.672 68.245 81.736 73.952 ;
      RECT 76.06 73.857 81.782 73.906 ;
      RECT 81.718 68.199 81.782 73.906 ;
      RECT 76.106 73.811 81.828 73.86 ;
      RECT 81.764 68.153 81.828 73.86 ;
      RECT 76.152 73.765 81.874 73.814 ;
      RECT 81.81 68.107 81.874 73.814 ;
      RECT 76.198 73.719 81.92 73.768 ;
      RECT 81.856 68.061 81.92 73.768 ;
      RECT 76.244 73.673 81.966 73.722 ;
      RECT 81.902 68.015 81.966 73.722 ;
      RECT 76.29 73.627 82.012 73.676 ;
      RECT 81.948 67.969 82.012 73.676 ;
      RECT 76.336 73.581 82.058 73.63 ;
      RECT 81.994 67.923 82.058 73.63 ;
      RECT 82.04 67.877 82.104 73.584 ;
      RECT 82.086 67.831 82.15 73.538 ;
      RECT 82.132 67.785 82.196 73.492 ;
      RECT 82.178 67.739 82.242 73.446 ;
      RECT 82.224 67.693 82.288 73.4 ;
      RECT 82.27 67.647 82.334 73.354 ;
      RECT 82.316 67.601 82.38 73.308 ;
      RECT 82.362 67.555 82.426 73.262 ;
      RECT 82.408 67.509 82.472 73.216 ;
      RECT 82.454 67.463 82.518 73.17 ;
      RECT 82.5 67.417 82.564 73.124 ;
      RECT 82.546 67.371 82.61 73.078 ;
      RECT 82.592 67.325 82.656 73.032 ;
      RECT 82.638 67.279 82.702 72.986 ;
      RECT 82.684 67.233 82.748 72.94 ;
      RECT 82.73 67.187 82.794 72.894 ;
      RECT 82.776 67.141 82.84 72.848 ;
      RECT 82.822 67.095 82.886 72.802 ;
      RECT 82.868 67.049 82.932 72.756 ;
      RECT 82.914 67.003 82.978 72.71 ;
      RECT 82.96 66.957 83.024 72.664 ;
      RECT 83.006 66.911 83.07 72.618 ;
      RECT 83.052 66.865 83.116 72.572 ;
      RECT 83.098 66.819 83.162 72.526 ;
      RECT 83.144 66.773 83.208 72.48 ;
      RECT 83.19 66.727 83.254 72.434 ;
      RECT 83.236 66.681 83.3 72.388 ;
      RECT 83.282 66.635 83.346 72.342 ;
      RECT 83.328 66.596 83.392 72.296 ;
      RECT 83.36 66.557 83.438 72.25 ;
      RECT 83.406 66.511 83.484 72.204 ;
      RECT 83.452 66.465 83.53 72.158 ;
      RECT 83.498 66.419 83.576 72.112 ;
      RECT 83.544 66.373 83.622 72.066 ;
      RECT 83.59 66.327 83.668 72.02 ;
      RECT 83.636 66.281 83.714 71.974 ;
      RECT 83.682 66.235 83.76 71.928 ;
      RECT 83.728 66.189 83.806 71.882 ;
      RECT 83.774 66.143 83.852 71.836 ;
      RECT 83.82 66.097 83.898 71.79 ;
      RECT 83.866 66.051 83.944 71.744 ;
      RECT 83.912 66.005 83.99 71.698 ;
      RECT 83.958 65.959 84.036 71.652 ;
      RECT 84.004 65.913 84.082 71.606 ;
      RECT 84.05 65.867 84.128 71.56 ;
      RECT 84.096 65.821 84.174 71.514 ;
      RECT 84.142 65.775 84.22 71.468 ;
      RECT 84.188 65.729 84.266 71.422 ;
      RECT 84.234 65.683 84.312 71.376 ;
      RECT 84.28 65.637 84.358 71.33 ;
      RECT 84.326 65.591 84.404 71.284 ;
      RECT 84.372 65.545 84.45 71.238 ;
      RECT 84.418 65.499 84.496 71.192 ;
      RECT 84.464 65.453 84.542 71.146 ;
      RECT 84.51 65.407 84.588 71.1 ;
      RECT 84.556 65.361 84.634 71.054 ;
      RECT 84.602 65.315 84.68 71.008 ;
      RECT 84.648 65.269 84.726 70.962 ;
      RECT 84.694 65.223 84.772 70.916 ;
      RECT 84.74 65.177 84.818 70.87 ;
      RECT 84.786 65.131 84.864 70.824 ;
      RECT 84.832 65.085 84.91 70.778 ;
      RECT 84.878 65.039 84.956 70.732 ;
      RECT 84.924 64.993 85.002 70.686 ;
      RECT 84.97 64.947 85.048 70.64 ;
      RECT 85.016 64.901 85.094 70.594 ;
      RECT 85.062 64.855 85.14 70.548 ;
      RECT 85.108 64.809 85.186 70.502 ;
      RECT 85.154 64.763 85.232 70.456 ;
      RECT 85.2 64.717 85.278 70.41 ;
      RECT 85.246 64.671 85.324 70.364 ;
      RECT 85.292 64.625 85.37 70.318 ;
      RECT 85.338 64.579 85.416 70.272 ;
      RECT 85.384 64.533 85.462 70.226 ;
      RECT 85.43 64.487 85.508 70.18 ;
      RECT 85.476 64.441 85.554 70.134 ;
      RECT 85.522 64.395 85.6 70.088 ;
      RECT 85.568 64.349 85.646 70.042 ;
      RECT 85.614 64.303 85.692 69.996 ;
      RECT 85.66 64.257 85.738 69.95 ;
      RECT 85.706 64.211 85.784 69.904 ;
      RECT 85.752 64.165 85.83 69.858 ;
      RECT 85.798 64.121 85.876 69.812 ;
      RECT 85.84 64.1 85.922 69.766 ;
      RECT 85.84 64.1 85.968 69.72 ;
      RECT 85.84 64.1 86.014 69.674 ;
      RECT 85.84 64.1 86.06 69.628 ;
      RECT 85.84 64.1 86.106 69.582 ;
      RECT 85.84 64.1 86.152 69.536 ;
      RECT 85.84 64.1 86.198 69.49 ;
      RECT 85.84 64.1 86.244 69.444 ;
      RECT 85.84 64.1 86.29 69.398 ;
      RECT 85.84 64.1 86.336 69.352 ;
      RECT 85.84 64.1 86.382 69.306 ;
      RECT 85.84 64.1 86.428 69.26 ;
      RECT 85.84 64.1 86.474 69.214 ;
      RECT 85.84 64.1 86.52 69.168 ;
      RECT 85.84 64.1 86.566 69.122 ;
      RECT 85.84 64.1 86.612 69.076 ;
      RECT 85.84 64.1 86.658 69.03 ;
      RECT 85.84 64.1 86.704 68.984 ;
      RECT 85.84 64.1 86.75 68.938 ;
      RECT 85.84 64.1 86.796 68.892 ;
      RECT 85.84 64.1 86.842 68.846 ;
      RECT 85.84 64.1 86.888 68.8 ;
      RECT 85.84 64.1 86.934 68.754 ;
      RECT 85.84 64.1 86.98 68.708 ;
      RECT 85.84 64.1 87.026 68.662 ;
      RECT 85.84 64.1 87.072 68.616 ;
      RECT 85.84 64.1 87.118 68.57 ;
      RECT 85.84 64.1 87.164 68.524 ;
      RECT 85.84 64.1 87.21 68.478 ;
      RECT 85.84 64.1 87.256 68.432 ;
      RECT 85.84 64.1 87.302 68.386 ;
      RECT 85.84 64.1 87.348 68.34 ;
      RECT 85.84 64.1 87.394 68.294 ;
      RECT 85.84 64.1 87.44 68.248 ;
      RECT 85.84 64.1 87.486 68.202 ;
      RECT 85.84 64.1 87.532 68.156 ;
      RECT 85.84 64.1 87.578 68.11 ;
      RECT 85.84 64.1 87.624 68.064 ;
      RECT 85.84 64.1 87.67 68.018 ;
      RECT 85.84 64.1 87.716 67.972 ;
      RECT 85.84 64.1 87.762 67.926 ;
      RECT 82.04 67.877 87.765 67.901 ;
      RECT 85.84 64.1 110 67.9 ;
      RECT 108.1 109.327 110 110 ;
      RECT 109.35 108.1 110 110 ;
      RECT 108.146 109.281 110 110 ;
      RECT 109.342 108.104 110 110 ;
      RECT 108.192 109.235 110 110 ;
      RECT 109.296 108.131 110 110 ;
      RECT 108.238 109.189 110 110 ;
      RECT 109.25 108.177 110 110 ;
      RECT 108.284 109.143 110 110 ;
      RECT 109.204 108.223 110 110 ;
      RECT 108.33 109.097 110 110 ;
      RECT 109.158 108.269 110 110 ;
      RECT 108.376 109.051 110 110 ;
      RECT 109.112 108.315 110 110 ;
      RECT 108.422 109.005 110 110 ;
      RECT 109.066 108.361 110 110 ;
      RECT 108.468 108.959 110 110 ;
      RECT 109.02 108.407 110 110 ;
      RECT 108.514 108.913 110 110 ;
      RECT 108.974 108.453 110 110 ;
      RECT 108.56 108.867 110 110 ;
      RECT 108.928 108.499 110 110 ;
      RECT 108.606 108.821 110 110 ;
      RECT 108.882 108.545 110 110 ;
      RECT 108.652 108.775 110 110 ;
      RECT 108.836 108.591 110 110 ;
      RECT 108.698 108.729 110 110 ;
      RECT 108.79 108.637 110 110 ;
      RECT 108.744 108.683 110 110 ;
      RECT 90.1 97.597 90.538 98.835 ;
      RECT 90.1 97.597 90.584 98.789 ;
      RECT 90.1 97.597 90.63 98.743 ;
      RECT 90.1 97.597 90.676 98.697 ;
      RECT 90.1 97.597 90.722 98.651 ;
      RECT 90.1 97.597 90.768 98.605 ;
      RECT 90.1 97.597 90.814 98.559 ;
      RECT 90.1 97.597 90.86 98.513 ;
      RECT 90.1 97.597 90.906 98.467 ;
      RECT 90.1 97.597 90.952 98.421 ;
      RECT 90.1 97.597 90.998 98.375 ;
      RECT 90.1 97.597 91.044 98.329 ;
      RECT 90.1 97.597 91.09 98.283 ;
      RECT 90.1 97.597 91.136 98.237 ;
      RECT 90.1 97.597 91.182 98.191 ;
      RECT 90.1 97.597 91.228 98.145 ;
      RECT 90.1 97.597 91.274 98.099 ;
      RECT 90.1 97.597 91.32 98.053 ;
      RECT 90.1 97.597 91.366 98.007 ;
      RECT 90.1 97.597 91.412 97.961 ;
      RECT 90.1 97.597 91.458 97.915 ;
      RECT 90.1 97.597 91.504 97.869 ;
      RECT 90.1 97.597 91.55 97.823 ;
      RECT 90.1 97.597 91.596 97.777 ;
      RECT 90.1 97.597 91.642 97.731 ;
      RECT 90.1 97.597 91.688 97.685 ;
      RECT 90.146 97.551 91.734 97.639 ;
      RECT 91.664 96.033 91.734 97.639 ;
      RECT 90.192 97.505 91.78 97.593 ;
      RECT 91.71 95.987 91.78 97.593 ;
      RECT 90.238 97.459 91.826 97.547 ;
      RECT 91.756 95.941 91.826 97.547 ;
      RECT 90.284 97.413 91.872 97.501 ;
      RECT 91.802 95.895 91.872 97.501 ;
      RECT 90.33 97.367 91.918 97.455 ;
      RECT 91.848 95.849 91.918 97.455 ;
      RECT 90.376 97.321 91.964 97.409 ;
      RECT 91.894 95.803 91.964 97.409 ;
      RECT 90.422 97.275 92.01 97.363 ;
      RECT 91.94 95.757 92.01 97.363 ;
      RECT 90.468 97.229 92.056 97.317 ;
      RECT 91.986 95.711 92.056 97.317 ;
      RECT 90.514 97.183 92.102 97.271 ;
      RECT 92.032 95.665 92.102 97.271 ;
      RECT 90.56 97.137 92.148 97.225 ;
      RECT 92.078 95.619 92.148 97.225 ;
      RECT 90.606 97.091 92.194 97.179 ;
      RECT 92.124 95.573 92.194 97.179 ;
      RECT 90.652 97.045 92.24 97.133 ;
      RECT 92.17 95.527 92.24 97.133 ;
      RECT 90.698 96.999 92.286 97.087 ;
      RECT 92.216 95.481 92.286 97.087 ;
      RECT 90.744 96.953 92.332 97.041 ;
      RECT 92.262 95.435 92.332 97.041 ;
      RECT 90.79 96.907 92.378 96.995 ;
      RECT 92.308 95.389 92.378 96.995 ;
      RECT 90.836 96.861 92.424 96.949 ;
      RECT 92.354 95.343 92.424 96.949 ;
      RECT 90.882 96.815 92.47 96.903 ;
      RECT 92.4 95.297 92.47 96.903 ;
      RECT 90.928 96.769 92.516 96.857 ;
      RECT 92.446 95.251 92.516 96.857 ;
      RECT 90.974 96.723 92.562 96.811 ;
      RECT 92.492 95.205 92.562 96.811 ;
      RECT 91.02 96.677 92.608 96.765 ;
      RECT 92.538 95.159 92.608 96.765 ;
      RECT 91.066 96.631 92.654 96.719 ;
      RECT 92.584 95.113 92.654 96.719 ;
      RECT 91.112 96.585 92.7 96.673 ;
      RECT 92.63 95.067 92.7 96.673 ;
      RECT 91.158 96.539 92.746 96.627 ;
      RECT 92.676 95.021 92.746 96.627 ;
      RECT 91.204 96.493 92.792 96.581 ;
      RECT 92.722 94.975 92.792 96.581 ;
      RECT 91.25 96.447 92.838 96.535 ;
      RECT 92.768 94.929 92.838 96.535 ;
      RECT 91.296 96.401 92.884 96.489 ;
      RECT 92.814 94.883 92.884 96.489 ;
      RECT 91.342 96.355 92.93 96.443 ;
      RECT 92.86 94.837 92.93 96.443 ;
      RECT 91.388 96.309 92.976 96.397 ;
      RECT 92.906 94.791 92.976 96.397 ;
      RECT 91.434 96.263 93.022 96.351 ;
      RECT 92.952 94.745 93.022 96.351 ;
      RECT 91.48 96.217 93.068 96.305 ;
      RECT 92.998 94.699 93.068 96.305 ;
      RECT 91.526 96.171 93.114 96.259 ;
      RECT 93.044 94.663 93.114 96.259 ;
      RECT 91.572 96.125 93.16 96.213 ;
      RECT 93.07 94.627 93.16 96.213 ;
      RECT 91.618 96.079 93.206 96.167 ;
      RECT 93.116 94.581 93.206 96.167 ;
      RECT 93.162 94.535 93.252 96.121 ;
      RECT 93.208 94.489 93.298 96.075 ;
      RECT 93.254 94.443 93.344 96.029 ;
      RECT 93.3 94.397 93.39 95.983 ;
      RECT 93.346 94.351 93.436 95.937 ;
      RECT 93.392 94.305 93.482 95.891 ;
      RECT 93.438 94.259 93.528 95.845 ;
      RECT 93.484 94.213 93.574 95.799 ;
      RECT 93.53 94.167 93.62 95.753 ;
      RECT 93.576 94.121 93.666 95.707 ;
      RECT 93.622 94.075 93.712 95.661 ;
      RECT 93.668 94.029 93.758 95.615 ;
      RECT 93.714 93.983 93.804 95.569 ;
      RECT 93.76 93.937 93.85 95.523 ;
      RECT 93.806 93.891 93.896 95.477 ;
      RECT 93.852 93.845 93.942 95.431 ;
      RECT 93.898 93.799 93.988 95.385 ;
      RECT 93.944 93.753 94.034 95.339 ;
      RECT 93.99 93.707 94.08 95.293 ;
      RECT 94.036 93.661 94.126 95.247 ;
      RECT 94.082 93.615 94.172 95.201 ;
      RECT 94.128 93.569 94.218 95.155 ;
      RECT 94.174 93.523 94.264 95.109 ;
      RECT 94.22 93.477 94.31 95.063 ;
      RECT 94.266 93.431 94.356 95.017 ;
      RECT 94.312 93.385 94.402 94.971 ;
      RECT 94.358 93.339 94.448 94.925 ;
      RECT 94.404 93.293 94.494 94.879 ;
      RECT 94.45 93.247 94.54 94.833 ;
      RECT 94.496 93.201 94.586 94.787 ;
      RECT 94.542 93.155 94.632 94.741 ;
      RECT 94.588 93.109 94.678 94.695 ;
      RECT 94.634 93.063 94.724 94.649 ;
      RECT 94.68 93.017 94.77 94.603 ;
      RECT 94.726 92.971 94.816 94.557 ;
      RECT 94.772 92.925 94.862 94.511 ;
      RECT 94.818 92.879 94.908 94.465 ;
      RECT 94.864 92.833 94.954 94.419 ;
      RECT 94.91 92.787 95 94.373 ;
      RECT 94.956 92.741 95.046 94.327 ;
      RECT 95.002 92.695 95.092 94.281 ;
      RECT 95.048 92.649 95.138 94.235 ;
      RECT 95.094 92.603 95.184 94.189 ;
      RECT 95.14 92.557 95.23 94.143 ;
      RECT 95.186 92.511 95.276 94.097 ;
      RECT 95.232 92.465 95.322 94.051 ;
      RECT 95.278 92.419 95.368 94.005 ;
      RECT 95.324 92.373 95.414 93.959 ;
      RECT 95.37 92.327 95.46 93.913 ;
      RECT 95.416 92.281 95.506 93.867 ;
      RECT 95.462 92.235 95.552 93.821 ;
      RECT 95.508 92.189 95.598 93.775 ;
      RECT 95.554 92.143 95.644 93.729 ;
      RECT 95.6 92.097 95.69 93.683 ;
      RECT 95.646 92.051 95.736 93.637 ;
      RECT 95.692 92.005 95.782 93.591 ;
      RECT 95.738 91.959 95.828 93.545 ;
      RECT 95.784 91.913 95.874 93.499 ;
      RECT 95.83 91.867 95.92 93.453 ;
      RECT 95.876 91.821 95.966 93.407 ;
      RECT 95.922 91.775 96.012 93.361 ;
      RECT 95.968 91.729 96.058 93.315 ;
      RECT 96.014 91.683 96.104 93.269 ;
      RECT 96.06 91.637 96.15 93.223 ;
      RECT 96.106 91.591 96.196 93.177 ;
      RECT 96.152 91.545 96.242 93.131 ;
      RECT 96.198 91.499 96.288 93.085 ;
      RECT 96.244 91.453 96.334 93.039 ;
      RECT 96.29 91.407 96.38 92.993 ;
      RECT 96.336 91.361 96.426 92.947 ;
      RECT 96.382 91.315 96.472 92.901 ;
      RECT 96.428 91.269 96.518 92.855 ;
      RECT 96.474 91.223 96.564 92.809 ;
      RECT 96.52 91.177 96.61 92.763 ;
      RECT 96.566 91.131 96.656 92.717 ;
      RECT 96.612 91.085 96.702 92.671 ;
      RECT 96.658 91.039 96.748 92.625 ;
      RECT 96.704 90.993 96.794 92.579 ;
      RECT 96.75 90.947 96.84 92.533 ;
      RECT 96.796 90.901 96.886 92.487 ;
      RECT 96.842 90.855 96.932 92.441 ;
      RECT 96.888 90.809 96.978 92.395 ;
      RECT 96.934 90.763 97.024 92.349 ;
      RECT 96.98 90.717 97.07 92.303 ;
      RECT 97.026 90.671 97.116 92.257 ;
      RECT 97.072 90.625 97.162 92.211 ;
      RECT 97.118 90.579 97.208 92.165 ;
      RECT 97.164 90.533 97.254 92.119 ;
      RECT 97.21 90.487 97.3 92.073 ;
      RECT 97.256 90.441 97.346 92.027 ;
      RECT 97.302 90.395 97.392 91.981 ;
      RECT 97.394 90.303 97.446 91.927 ;
      RECT 97.44 90.257 97.492 91.881 ;
      RECT 97.486 90.211 97.538 91.835 ;
      RECT 97.532 90.165 97.584 91.789 ;
      RECT 97.578 90.121 97.63 91.743 ;
      RECT 97.62 90.1 97.676 91.697 ;
      RECT 97.348 90.349 97.4 91.954 ;
      RECT 97.62 90.1 97.722 91.651 ;
      RECT 97.62 90.1 97.768 91.605 ;
      RECT 97.62 90.1 97.814 91.559 ;
      RECT 97.62 90.1 97.86 91.513 ;
      RECT 97.62 90.1 97.906 91.467 ;
      RECT 97.62 90.1 97.952 91.421 ;
      RECT 97.62 90.1 97.998 91.375 ;
      RECT 97.62 90.1 98.044 91.329 ;
      RECT 97.62 90.1 98.09 91.283 ;
      RECT 97.62 90.1 98.136 91.237 ;
      RECT 97.62 90.1 98.182 91.191 ;
      RECT 97.62 90.1 98.228 91.145 ;
      RECT 97.62 90.1 98.274 91.099 ;
      RECT 97.62 90.1 98.32 91.053 ;
      RECT 97.62 90.1 98.366 91.007 ;
      RECT 97.62 90.1 98.412 90.961 ;
      RECT 97.62 90.1 98.458 90.915 ;
      RECT 97.62 90.1 98.504 90.869 ;
      RECT 97.62 90.1 98.55 90.823 ;
      RECT 97.62 90.1 98.596 90.777 ;
      RECT 97.62 90.1 98.642 90.731 ;
      RECT 97.62 90.1 98.688 90.685 ;
      RECT 97.62 90.1 98.734 90.639 ;
      RECT 97.62 90.1 98.78 90.593 ;
      RECT 97.62 90.1 98.826 90.547 ;
      RECT 97.62 90.1 98.872 90.501 ;
      RECT 43.1 75.057 43.538 75.55 ;
      RECT 43.1 75.057 43.584 75.504 ;
      RECT 43.1 75.057 43.63 75.458 ;
      RECT 43.1 75.057 43.676 75.412 ;
      RECT 43.1 75.057 43.722 75.366 ;
      RECT 43.1 75.057 43.768 75.32 ;
      RECT 43.1 75.057 43.814 75.274 ;
      RECT 43.1 75.057 43.86 75.228 ;
      RECT 43.1 75.057 43.906 75.182 ;
      RECT 43.1 75.057 43.952 75.136 ;
      RECT 43.146 75.011 43.998 75.09 ;
      RECT 43.192 74.965 44.044 75.044 ;
      RECT 43.238 74.919 44.09 74.998 ;
      RECT 43.284 74.873 44.136 74.952 ;
      RECT 43.33 74.827 44.182 74.906 ;
      RECT 43.376 74.781 44.228 74.86 ;
      RECT 43.422 74.735 44.274 74.814 ;
      RECT 43.468 74.689 44.32 74.768 ;
      RECT 43.514 74.643 44.366 74.722 ;
      RECT 43.56 74.597 44.412 74.676 ;
      RECT 43.606 74.551 44.458 74.63 ;
      RECT 43.652 74.505 44.504 74.584 ;
      RECT 43.698 74.459 44.55 74.538 ;
      RECT 43.744 74.413 44.596 74.492 ;
      RECT 43.79 74.367 44.642 74.446 ;
      RECT 43.836 74.321 44.688 74.4 ;
      RECT 43.882 74.275 44.734 74.354 ;
      RECT 43.928 74.229 44.78 74.308 ;
      RECT 43.974 74.183 44.826 74.262 ;
      RECT 44.02 74.137 44.872 74.216 ;
      RECT 44.066 74.091 44.918 74.17 ;
      RECT 44.112 74.045 44.964 74.124 ;
      RECT 44.158 73.999 45.01 74.078 ;
      RECT 44.204 73.953 45.056 74.032 ;
      RECT 44.25 73.907 45.102 73.986 ;
      RECT 44.296 73.861 45.148 73.94 ;
      RECT 44.342 73.815 45.194 73.894 ;
      RECT 44.388 73.769 45.24 73.848 ;
      RECT 44.434 73.723 45.286 73.802 ;
      RECT 44.48 73.677 45.332 73.756 ;
      RECT 44.526 73.631 45.378 73.71 ;
      RECT 44.572 73.585 45.424 73.664 ;
      RECT 44.618 73.539 45.47 73.618 ;
      RECT 44.664 73.493 45.516 73.572 ;
      RECT 44.71 73.447 45.562 73.526 ;
      RECT 44.756 73.401 45.608 73.48 ;
      RECT 44.802 73.355 45.654 73.434 ;
      RECT 44.848 73.309 45.7 73.388 ;
      RECT 44.894 73.263 45.746 73.342 ;
      RECT 44.94 73.217 45.792 73.296 ;
      RECT 44.986 73.171 45.838 73.25 ;
      RECT 45.032 73.125 45.884 73.204 ;
      RECT 45.078 73.079 45.93 73.158 ;
      RECT 45.124 73.033 45.976 73.112 ;
      RECT 45.17 72.987 46.022 73.066 ;
      RECT 45.216 72.941 46.068 73.02 ;
      RECT 45.262 72.895 46.114 72.974 ;
      RECT 45.308 72.849 46.16 72.928 ;
      RECT 45.354 72.803 46.206 72.882 ;
      RECT 45.4 72.757 46.252 72.836 ;
      RECT 45.446 72.711 46.298 72.79 ;
      RECT 45.492 72.665 46.344 72.744 ;
      RECT 45.538 72.619 46.39 72.698 ;
      RECT 45.584 72.573 46.436 72.652 ;
      RECT 45.63 72.527 46.482 72.606 ;
      RECT 45.676 72.481 46.528 72.56 ;
      RECT 45.722 72.435 46.574 72.514 ;
      RECT 45.768 72.389 46.62 72.468 ;
      RECT 45.814 72.343 46.666 72.422 ;
      RECT 45.86 72.297 46.712 72.376 ;
      RECT 45.906 72.251 46.758 72.33 ;
      RECT 45.952 72.205 46.804 72.284 ;
      RECT 45.998 72.159 46.85 72.238 ;
      RECT 46.044 72.113 46.896 72.192 ;
      RECT 46.09 72.067 46.942 72.146 ;
      RECT 46.136 72.021 46.988 72.1 ;
      RECT 46.182 71.975 47.034 72.054 ;
      RECT 46.228 71.929 47.08 72.008 ;
      RECT 46.274 71.883 47.126 71.962 ;
      RECT 46.32 71.837 47.172 71.916 ;
      RECT 46.366 71.791 47.218 71.87 ;
      RECT 46.412 71.745 47.264 71.824 ;
      RECT 46.458 71.699 47.31 71.778 ;
      RECT 46.504 71.653 47.356 71.732 ;
      RECT 46.55 71.607 47.402 71.686 ;
      RECT 46.596 71.561 47.448 71.64 ;
      RECT 46.642 71.515 47.494 71.594 ;
      RECT 46.688 71.469 47.54 71.548 ;
      RECT 46.734 71.423 47.586 71.502 ;
      RECT 46.78 71.377 47.632 71.456 ;
      RECT 46.826 71.331 47.678 71.41 ;
      RECT 46.872 71.285 47.724 71.364 ;
      RECT 46.918 71.239 47.77 71.318 ;
      RECT 46.964 71.193 47.816 71.272 ;
      RECT 47.01 71.147 47.862 71.226 ;
      RECT 47.056 71.101 47.908 71.18 ;
      RECT 47.102 71.055 47.954 71.134 ;
      RECT 47.148 71.009 48 71.088 ;
      RECT 47.194 70.963 48.046 71.042 ;
      RECT 47.24 70.917 48.092 70.996 ;
      RECT 47.286 70.871 48.138 70.95 ;
      RECT 47.332 70.825 48.184 70.904 ;
      RECT 47.378 70.779 48.23 70.858 ;
      RECT 47.424 70.733 48.276 70.812 ;
      RECT 47.47 70.687 48.322 70.766 ;
      RECT 47.516 70.641 48.368 70.72 ;
      RECT 47.562 70.595 48.414 70.674 ;
      RECT 47.608 70.549 48.46 70.628 ;
      RECT 47.654 70.503 48.506 70.582 ;
      RECT 47.7 70.457 48.552 70.536 ;
      RECT 47.746 70.411 48.598 70.49 ;
      RECT 47.792 70.365 48.644 70.444 ;
      RECT 47.838 70.319 48.69 70.398 ;
      RECT 47.884 70.273 48.736 70.352 ;
      RECT 47.93 70.227 48.782 70.306 ;
      RECT 47.976 70.181 48.828 70.26 ;
      RECT 48.022 70.135 48.874 70.214 ;
      RECT 48.068 70.089 48.92 70.168 ;
      RECT 48.114 70.043 48.966 70.122 ;
      RECT 48.16 69.997 49.012 70.076 ;
      RECT 48.206 69.951 49.058 70.03 ;
      RECT 48.252 69.905 49.104 69.984 ;
      RECT 48.298 69.859 49.15 69.938 ;
      RECT 48.344 69.813 49.196 69.892 ;
      RECT 48.39 69.767 49.242 69.846 ;
      RECT 48.436 69.721 49.288 69.8 ;
      RECT 48.482 69.675 49.334 69.754 ;
      RECT 48.528 69.629 49.38 69.708 ;
      RECT 48.574 69.583 49.426 69.662 ;
      RECT 48.62 69.537 49.472 69.616 ;
      RECT 48.666 69.491 49.518 69.57 ;
      RECT 48.712 69.445 49.564 69.524 ;
      RECT 48.758 69.399 49.61 69.478 ;
      RECT 48.804 69.353 49.656 69.432 ;
      RECT 48.85 69.307 49.702 69.386 ;
      RECT 48.896 69.261 49.748 69.34 ;
      RECT 48.942 69.215 49.794 69.294 ;
      RECT 48.988 69.169 49.84 69.248 ;
      RECT 49.034 69.123 49.886 69.202 ;
      RECT 49.08 69.077 49.932 69.156 ;
      RECT 49.126 69.031 49.978 69.11 ;
      RECT 49.172 68.985 50.024 69.064 ;
      RECT 49.218 68.939 50.07 69.018 ;
      RECT 49.264 68.893 50.116 68.972 ;
      RECT 49.31 68.847 50.162 68.926 ;
      RECT 49.356 68.801 50.208 68.88 ;
      RECT 49.402 68.755 50.254 68.834 ;
      RECT 49.448 68.709 50.3 68.788 ;
      RECT 49.494 68.663 50.346 68.742 ;
      RECT 49.54 68.617 50.392 68.696 ;
      RECT 49.586 68.571 50.438 68.65 ;
      RECT 49.632 68.525 50.484 68.604 ;
      RECT 49.678 68.479 50.53 68.558 ;
      RECT 49.724 68.433 50.576 68.512 ;
      RECT 49.77 68.387 50.622 68.466 ;
      RECT 49.816 68.341 50.668 68.42 ;
      RECT 49.862 68.295 50.714 68.374 ;
      RECT 49.908 68.249 50.76 68.328 ;
      RECT 49.954 68.203 50.806 68.282 ;
      RECT 50 68.157 50.852 68.236 ;
      RECT 50.046 68.111 50.898 68.19 ;
      RECT 50.092 68.065 50.944 68.144 ;
      RECT 50.138 68.019 50.99 68.098 ;
      RECT 50.184 67.973 51.036 68.052 ;
      RECT 50.23 67.927 51.082 68.006 ;
      RECT 50.276 67.881 51.128 67.96 ;
      RECT 50.322 67.835 51.174 67.914 ;
      RECT 50.368 67.789 51.22 67.868 ;
      RECT 50.414 67.743 51.266 67.822 ;
      RECT 50.46 67.697 51.312 67.776 ;
      RECT 50.506 67.651 51.358 67.73 ;
      RECT 50.552 67.605 51.404 67.684 ;
      RECT 50.598 67.559 51.45 67.638 ;
      RECT 50.644 67.513 51.496 67.592 ;
      RECT 50.69 67.467 51.542 67.546 ;
      RECT 50.736 67.421 51.588 67.5 ;
      RECT 50.782 67.375 51.634 67.454 ;
      RECT 50.828 67.329 51.68 67.408 ;
      RECT 50.874 67.283 51.726 67.362 ;
      RECT 50.92 67.237 51.772 67.316 ;
      RECT 50.966 67.191 51.818 67.27 ;
      RECT 51.012 67.145 51.864 67.224 ;
      RECT 51.058 67.099 51.91 67.178 ;
      RECT 51.104 67.053 51.956 67.132 ;
      RECT 51.15 67.007 52.002 67.086 ;
      RECT 51.196 66.961 52.048 67.04 ;
      RECT 51.242 66.915 52.094 66.994 ;
      RECT 51.288 66.869 52.14 66.948 ;
      RECT 51.334 66.823 52.186 66.902 ;
      RECT 51.38 66.777 52.232 66.856 ;
      RECT 51.426 66.731 52.278 66.81 ;
      RECT 51.472 66.685 52.324 66.764 ;
      RECT 51.518 66.639 52.37 66.718 ;
      RECT 51.564 66.593 52.416 66.672 ;
      RECT 51.61 66.547 52.462 66.626 ;
      RECT 51.656 66.501 52.508 66.58 ;
      RECT 51.702 66.455 52.554 66.534 ;
      RECT 51.748 66.409 52.6 66.488 ;
      RECT 51.794 66.363 52.646 66.442 ;
      RECT 51.84 66.317 52.692 66.396 ;
      RECT 51.886 66.271 52.738 66.35 ;
      RECT 51.932 66.225 52.784 66.304 ;
      RECT 51.978 66.179 52.83 66.258 ;
      RECT 52.024 66.133 52.876 66.212 ;
      RECT 52.07 66.087 52.922 66.166 ;
      RECT 52.116 66.041 52.968 66.12 ;
      RECT 52.162 65.995 53.014 66.074 ;
      RECT 52.208 65.949 53.06 66.028 ;
      RECT 52.254 65.903 53.106 65.982 ;
      RECT 52.3 65.857 53.152 65.936 ;
      RECT 52.346 65.811 53.198 65.89 ;
      RECT 52.392 65.765 53.244 65.844 ;
      RECT 52.438 65.719 53.29 65.798 ;
      RECT 52.484 65.673 53.336 65.752 ;
      RECT 52.53 65.627 53.382 65.706 ;
      RECT 52.576 65.581 53.428 65.66 ;
      RECT 52.622 65.535 53.474 65.614 ;
      RECT 52.668 65.489 53.52 65.568 ;
      RECT 52.714 65.443 53.566 65.522 ;
      RECT 52.76 65.397 53.612 65.476 ;
      RECT 52.806 65.351 53.658 65.43 ;
      RECT 52.852 65.305 53.704 65.384 ;
      RECT 52.898 65.259 53.75 65.338 ;
      RECT 52.944 65.213 53.796 65.292 ;
      RECT 52.99 65.167 53.842 65.246 ;
      RECT 53.036 65.121 53.888 65.2 ;
      RECT 53.082 65.075 53.934 65.154 ;
      RECT 53.128 65.029 53.98 65.108 ;
      RECT 53.174 64.983 54.026 65.062 ;
      RECT 53.22 64.937 54.072 65.016 ;
      RECT 53.266 64.891 54.118 64.97 ;
      RECT 53.312 64.845 54.164 64.924 ;
      RECT 53.358 64.799 54.21 64.878 ;
      RECT 53.404 64.753 54.256 64.832 ;
      RECT 53.45 64.707 54.302 64.786 ;
      RECT 53.496 64.661 54.348 64.74 ;
      RECT 53.542 64.615 54.394 64.694 ;
      RECT 53.588 64.569 54.44 64.648 ;
      RECT 53.634 64.523 54.486 64.602 ;
      RECT 53.68 64.477 54.532 64.556 ;
      RECT 53.726 64.431 54.578 64.51 ;
      RECT 53.772 64.385 54.624 64.464 ;
      RECT 53.818 64.339 54.67 64.418 ;
      RECT 53.864 64.293 54.716 64.372 ;
      RECT 53.91 64.247 54.762 64.326 ;
      RECT 53.956 64.201 54.808 64.28 ;
      RECT 54.002 64.155 54.854 64.234 ;
      RECT 54.048 64.109 54.9 64.188 ;
      RECT 54.094 64.063 54.946 64.142 ;
      RECT 54.14 64.017 54.992 64.096 ;
      RECT 54.186 63.971 55.038 64.05 ;
      RECT 54.232 63.925 55.084 64.004 ;
      RECT 54.278 63.879 55.13 63.958 ;
      RECT 54.324 63.833 55.176 63.912 ;
      RECT 54.37 63.787 55.222 63.866 ;
      RECT 54.416 63.741 55.268 63.82 ;
      RECT 54.462 63.695 55.314 63.774 ;
      RECT 54.508 63.649 55.36 63.728 ;
      RECT 54.554 63.603 55.4 63.685 ;
      RECT 54.6 63.557 55.446 63.642 ;
      RECT 54.646 63.511 55.492 63.596 ;
      RECT 54.692 63.465 55.538 63.55 ;
      RECT 54.738 63.419 55.584 63.504 ;
      RECT 54.784 63.373 55.63 63.458 ;
      RECT 54.83 63.327 55.676 63.412 ;
      RECT 54.876 63.281 55.722 63.366 ;
      RECT 54.922 63.235 55.768 63.32 ;
      RECT 54.968 63.189 55.814 63.274 ;
      RECT 55.014 63.143 55.86 63.228 ;
      RECT 55.06 63.097 55.906 63.182 ;
      RECT 55.106 63.051 55.952 63.136 ;
      RECT 55.152 63.005 55.998 63.09 ;
      RECT 55.198 62.959 56.044 63.044 ;
      RECT 55.244 62.913 56.09 62.998 ;
      RECT 55.29 62.867 56.136 62.952 ;
      RECT 55.336 62.821 56.182 62.906 ;
      RECT 55.382 62.775 56.228 62.86 ;
      RECT 55.428 62.729 56.274 62.814 ;
      RECT 55.474 62.683 56.32 62.768 ;
      RECT 55.52 62.637 56.366 62.722 ;
      RECT 55.566 62.591 56.412 62.676 ;
      RECT 55.612 62.545 56.458 62.63 ;
      RECT 55.658 62.499 56.504 62.584 ;
      RECT 55.704 62.453 56.55 62.538 ;
      RECT 55.75 62.407 56.596 62.492 ;
      RECT 55.796 62.361 56.642 62.446 ;
      RECT 55.842 62.315 56.688 62.4 ;
      RECT 55.888 62.269 56.734 62.354 ;
      RECT 55.934 62.223 56.78 62.308 ;
      RECT 55.98 62.177 56.826 62.262 ;
      RECT 56.026 62.131 56.872 62.216 ;
      RECT 56.072 62.085 56.918 62.17 ;
      RECT 56.118 62.039 56.964 62.124 ;
      RECT 56.164 61.993 57.01 62.078 ;
      RECT 56.21 61.947 57.056 62.032 ;
      RECT 56.256 61.901 57.102 61.986 ;
      RECT 56.302 61.855 57.148 61.94 ;
      RECT 56.348 61.809 57.194 61.894 ;
      RECT 56.394 61.763 57.24 61.848 ;
      RECT 56.44 61.717 57.286 61.802 ;
      RECT 56.486 61.671 57.332 61.756 ;
      RECT 56.532 61.625 57.378 61.71 ;
      RECT 56.578 61.579 57.424 61.664 ;
      RECT 56.624 61.533 57.47 61.618 ;
      RECT 56.67 61.487 57.516 61.572 ;
      RECT 56.716 61.441 57.562 61.526 ;
      RECT 56.762 61.395 57.608 61.48 ;
      RECT 56.808 61.349 57.654 61.434 ;
      RECT 56.854 61.303 57.7 61.388 ;
      RECT 56.9 61.257 57.746 61.342 ;
      RECT 56.946 61.211 57.792 61.296 ;
      RECT 56.992 61.165 57.838 61.25 ;
      RECT 57.038 61.119 57.884 61.204 ;
      RECT 57.084 61.073 57.93 61.158 ;
      RECT 57.13 61.027 57.976 61.112 ;
      RECT 57.176 60.981 58.022 61.066 ;
      RECT 57.222 60.935 58.068 61.02 ;
      RECT 57.268 60.889 58.114 60.974 ;
      RECT 57.314 60.843 58.16 60.928 ;
      RECT 57.36 60.797 58.206 60.882 ;
      RECT 57.406 60.751 58.252 60.836 ;
      RECT 57.452 60.705 58.298 60.79 ;
      RECT 57.498 60.659 58.344 60.744 ;
      RECT 57.544 60.613 58.39 60.698 ;
      RECT 57.59 60.567 58.436 60.652 ;
      RECT 57.636 60.521 58.482 60.606 ;
      RECT 57.682 60.475 58.528 60.56 ;
      RECT 57.728 60.429 58.574 60.514 ;
      RECT 57.774 60.383 58.62 60.468 ;
      RECT 57.82 60.337 58.666 60.422 ;
      RECT 57.866 60.291 58.712 60.376 ;
      RECT 57.912 60.245 58.758 60.33 ;
      RECT 57.958 60.199 58.804 60.284 ;
      RECT 58.004 60.153 58.85 60.238 ;
      RECT 58.05 60.107 58.896 60.192 ;
      RECT 58.096 60.061 58.942 60.146 ;
      RECT 58.142 60.015 58.988 60.1 ;
      RECT 58.188 59.969 59.034 60.054 ;
      RECT 58.234 59.923 59.08 60.008 ;
      RECT 58.28 59.877 59.126 59.962 ;
      RECT 58.326 59.831 59.172 59.916 ;
      RECT 58.372 59.785 59.218 59.87 ;
      RECT 58.418 59.739 59.264 59.824 ;
      RECT 58.464 59.693 59.31 59.778 ;
      RECT 58.51 59.647 59.356 59.732 ;
      RECT 58.556 59.601 59.402 59.686 ;
      RECT 58.602 59.555 59.448 59.64 ;
      RECT 58.648 59.509 59.494 59.594 ;
      RECT 58.694 59.463 59.54 59.548 ;
      RECT 58.74 59.417 59.586 59.502 ;
      RECT 58.786 59.371 59.632 59.456 ;
      RECT 58.832 59.325 59.678 59.41 ;
      RECT 58.878 59.279 59.724 59.364 ;
      RECT 58.924 59.233 59.77 59.318 ;
      RECT 58.97 59.187 59.816 59.272 ;
      RECT 59.016 59.141 59.862 59.226 ;
      RECT 59.062 59.095 59.908 59.18 ;
      RECT 59.108 59.049 59.954 59.134 ;
      RECT 59.154 59.003 60 59.088 ;
      RECT 59.2 58.957 60.046 59.042 ;
      RECT 59.246 58.911 60.092 58.996 ;
      RECT 59.292 58.865 60.138 58.95 ;
      RECT 59.338 58.819 60.184 58.904 ;
      RECT 59.384 58.773 60.23 58.858 ;
      RECT 59.43 58.727 60.276 58.812 ;
      RECT 59.476 58.681 60.322 58.766 ;
      RECT 59.522 58.635 60.368 58.72 ;
      RECT 59.568 58.589 60.414 58.674 ;
      RECT 59.614 58.543 60.46 58.628 ;
      RECT 59.66 58.497 60.506 58.582 ;
      RECT 59.706 58.451 60.552 58.536 ;
      RECT 59.752 58.405 60.598 58.49 ;
      RECT 59.798 58.359 60.644 58.444 ;
      RECT 59.844 58.313 60.69 58.398 ;
      RECT 59.89 58.267 60.736 58.352 ;
      RECT 59.936 58.221 60.782 58.306 ;
      RECT 59.982 58.175 60.828 58.26 ;
      RECT 60.028 58.129 60.874 58.214 ;
      RECT 60.074 58.083 60.92 58.168 ;
      RECT 60.12 58.037 60.966 58.122 ;
      RECT 60.166 57.991 61.012 58.076 ;
      RECT 60.212 57.945 61.058 58.03 ;
      RECT 60.258 57.899 61.104 57.984 ;
      RECT 60.304 57.853 61.15 57.938 ;
      RECT 60.35 57.807 61.196 57.892 ;
      RECT 60.396 57.761 61.242 57.846 ;
      RECT 60.442 57.715 61.288 57.8 ;
      RECT 60.488 57.669 61.334 57.754 ;
      RECT 60.534 57.623 61.38 57.708 ;
      RECT 60.58 57.577 61.426 57.662 ;
      RECT 60.626 57.531 61.472 57.616 ;
      RECT 60.672 57.485 61.518 57.57 ;
      RECT 60.718 57.439 61.564 57.524 ;
      RECT 60.764 57.393 61.61 57.478 ;
      RECT 60.81 57.347 61.656 57.432 ;
      RECT 60.856 57.301 61.702 57.386 ;
      RECT 60.902 57.255 61.748 57.34 ;
      RECT 60.948 57.209 61.794 57.294 ;
      RECT 60.994 57.163 61.84 57.248 ;
      RECT 61.04 57.117 61.886 57.202 ;
      RECT 61.086 57.071 61.932 57.156 ;
      RECT 61.132 57.025 61.978 57.11 ;
      RECT 61.178 56.979 62.024 57.064 ;
      RECT 61.224 56.933 62.07 57.018 ;
      RECT 61.27 56.887 62.116 56.972 ;
      RECT 61.316 56.841 62.162 56.926 ;
      RECT 61.362 56.795 62.208 56.88 ;
      RECT 61.408 56.749 62.254 56.834 ;
      RECT 61.454 56.703 62.3 56.788 ;
      RECT 61.5 56.657 62.346 56.742 ;
      RECT 61.546 56.611 62.392 56.696 ;
      RECT 61.592 56.565 62.438 56.65 ;
      RECT 61.638 56.519 62.484 56.604 ;
      RECT 61.684 56.473 62.53 56.558 ;
      RECT 61.73 56.427 62.576 56.512 ;
      RECT 61.776 56.381 62.622 56.466 ;
      RECT 61.822 56.335 62.668 56.42 ;
      RECT 61.868 56.289 62.714 56.374 ;
      RECT 61.914 56.243 62.76 56.328 ;
      RECT 61.96 56.197 62.806 56.282 ;
      RECT 62.006 56.151 62.852 56.236 ;
      RECT 62.052 56.105 62.898 56.19 ;
      RECT 62.098 56.059 62.944 56.144 ;
      RECT 62.144 56.013 62.99 56.098 ;
      RECT 62.19 55.967 63.036 56.052 ;
      RECT 62.236 55.921 63.082 56.006 ;
      RECT 62.282 55.875 63.128 55.96 ;
      RECT 62.328 55.829 63.174 55.914 ;
      RECT 62.374 55.783 63.22 55.868 ;
      RECT 62.42 55.737 63.266 55.822 ;
      RECT 62.466 55.691 63.312 55.776 ;
      RECT 62.512 55.645 63.358 55.73 ;
      RECT 62.558 55.599 63.404 55.684 ;
      RECT 62.604 55.553 63.45 55.638 ;
      RECT 62.65 55.507 63.496 55.592 ;
      RECT 62.696 55.461 63.542 55.546 ;
      RECT 62.742 55.415 63.588 55.5 ;
      RECT 62.788 55.369 63.634 55.454 ;
      RECT 62.834 55.323 63.68 55.408 ;
      RECT 62.88 55.277 63.726 55.362 ;
      RECT 62.926 55.231 63.772 55.316 ;
      RECT 62.972 55.185 63.818 55.27 ;
      RECT 63.018 55.139 63.864 55.224 ;
      RECT 63.064 55.093 63.91 55.178 ;
      RECT 63.11 55.047 63.956 55.132 ;
      RECT 63.156 55.001 64.002 55.086 ;
      RECT 63.202 54.955 64.048 55.04 ;
      RECT 63.248 54.909 64.094 54.994 ;
      RECT 63.294 54.863 64.14 54.948 ;
      RECT 63.34 54.817 64.186 54.902 ;
      RECT 63.386 54.771 64.232 54.856 ;
      RECT 63.432 54.725 64.278 54.81 ;
      RECT 63.478 54.679 64.324 54.764 ;
      RECT 63.524 54.633 64.37 54.718 ;
      RECT 63.57 54.587 64.416 54.672 ;
      RECT 63.616 54.541 64.462 54.626 ;
      RECT 63.662 54.495 64.508 54.58 ;
      RECT 63.708 54.449 64.554 54.534 ;
      RECT 63.754 54.403 64.6 54.488 ;
      RECT 63.8 54.357 64.646 54.442 ;
      RECT 63.846 54.311 64.692 54.396 ;
      RECT 63.892 54.265 64.738 54.35 ;
      RECT 63.938 54.219 64.784 54.304 ;
      RECT 63.984 54.173 64.83 54.258 ;
      RECT 64.03 54.127 64.876 54.212 ;
      RECT 64.076 54.081 64.922 54.166 ;
      RECT 64.122 54.035 64.968 54.12 ;
      RECT 64.168 53.989 65.014 54.074 ;
      RECT 64.214 53.943 65.06 54.028 ;
      RECT 64.26 53.897 65.106 53.982 ;
      RECT 64.306 53.851 65.152 53.936 ;
      RECT 64.352 53.805 65.198 53.89 ;
      RECT 64.398 53.759 65.244 53.844 ;
      RECT 64.444 53.713 65.29 53.798 ;
      RECT 64.49 53.667 65.336 53.752 ;
      RECT 64.536 53.621 65.382 53.706 ;
      RECT 64.582 53.575 65.428 53.66 ;
      RECT 64.628 53.529 65.474 53.614 ;
      RECT 64.674 53.483 65.52 53.568 ;
      RECT 64.72 53.437 65.566 53.522 ;
      RECT 64.766 53.391 65.612 53.476 ;
      RECT 64.812 53.345 65.658 53.43 ;
      RECT 64.858 53.299 65.704 53.384 ;
      RECT 64.904 53.253 65.75 53.338 ;
      RECT 64.95 53.207 65.796 53.292 ;
      RECT 64.996 53.161 65.842 53.246 ;
      RECT 65.042 53.115 65.888 53.2 ;
      RECT 65.088 53.069 65.934 53.154 ;
      RECT 65.134 53.023 65.98 53.108 ;
      RECT 65.18 52.977 66.026 53.062 ;
      RECT 65.226 52.931 66.072 53.016 ;
      RECT 65.272 52.885 66.118 52.97 ;
      RECT 65.318 52.839 66.164 52.924 ;
      RECT 65.364 52.793 66.21 52.878 ;
      RECT 65.41 52.747 66.256 52.832 ;
      RECT 65.456 52.701 66.302 52.786 ;
      RECT 65.502 52.655 66.348 52.74 ;
      RECT 65.548 52.609 66.394 52.694 ;
      RECT 65.594 52.563 66.44 52.648 ;
      RECT 65.64 52.517 66.486 52.602 ;
      RECT 65.686 52.471 66.532 52.556 ;
      RECT 65.732 52.425 66.578 52.51 ;
      RECT 65.778 52.379 66.624 52.464 ;
      RECT 65.824 52.333 66.67 52.418 ;
      RECT 65.87 52.287 66.716 52.372 ;
      RECT 65.916 52.241 66.762 52.326 ;
      RECT 65.962 52.195 66.808 52.28 ;
      RECT 66.008 52.149 66.854 52.234 ;
      RECT 66.054 52.103 66.9 52.188 ;
      RECT 66.1 52.057 66.946 52.142 ;
      RECT 66.146 52.011 66.992 52.096 ;
      RECT 66.192 51.965 67.038 52.05 ;
      RECT 66.238 51.919 67.084 52.004 ;
      RECT 66.284 51.873 67.13 51.958 ;
      RECT 66.33 51.827 67.176 51.912 ;
      RECT 66.376 51.781 67.222 51.866 ;
      RECT 66.422 51.735 67.268 51.82 ;
      RECT 66.468 51.689 67.314 51.774 ;
      RECT 66.514 51.643 67.36 51.728 ;
      RECT 66.56 51.597 67.406 51.682 ;
      RECT 66.606 51.551 67.452 51.636 ;
      RECT 66.652 51.505 67.498 51.59 ;
      RECT 66.698 51.459 67.544 51.544 ;
      RECT 66.744 51.413 67.59 51.498 ;
      RECT 66.79 51.367 67.636 51.452 ;
      RECT 66.836 51.321 67.682 51.406 ;
      RECT 66.882 51.275 67.728 51.36 ;
      RECT 66.928 51.229 67.774 51.314 ;
      RECT 66.974 51.183 67.82 51.268 ;
      RECT 67.02 51.137 67.866 51.222 ;
      RECT 67.066 51.091 67.912 51.176 ;
      RECT 67.112 51.045 67.958 51.13 ;
      RECT 67.158 50.999 68.004 51.084 ;
      RECT 67.204 50.953 68.05 51.038 ;
      RECT 67.25 50.907 68.096 50.992 ;
      RECT 67.296 50.861 68.142 50.946 ;
      RECT 67.342 50.815 68.188 50.9 ;
      RECT 67.388 50.769 68.234 50.854 ;
      RECT 67.434 50.723 68.28 50.808 ;
      RECT 67.48 50.677 68.326 50.762 ;
      RECT 67.526 50.631 68.372 50.716 ;
      RECT 67.572 50.585 68.418 50.67 ;
      RECT 67.618 50.539 68.464 50.624 ;
      RECT 67.664 50.493 68.51 50.578 ;
      RECT 67.71 50.447 68.556 50.532 ;
      RECT 67.756 50.401 68.602 50.486 ;
      RECT 67.802 50.355 68.648 50.44 ;
      RECT 67.848 50.309 68.694 50.394 ;
      RECT 67.894 50.263 68.74 50.348 ;
      RECT 67.94 50.217 68.786 50.302 ;
      RECT 67.986 50.171 68.832 50.256 ;
      RECT 68.032 50.125 68.878 50.21 ;
      RECT 68.078 50.079 68.924 50.164 ;
      RECT 68.124 50.033 68.97 50.118 ;
      RECT 68.17 49.987 69.016 50.072 ;
      RECT 68.216 49.941 69.062 50.026 ;
      RECT 68.262 49.895 69.108 49.98 ;
      RECT 68.308 49.849 69.154 49.934 ;
      RECT 68.354 49.803 69.2 49.888 ;
      RECT 68.4 49.757 69.246 49.842 ;
      RECT 68.446 49.711 69.292 49.796 ;
      RECT 68.492 49.665 69.338 49.75 ;
      RECT 68.538 49.619 69.384 49.704 ;
      RECT 68.584 49.573 69.43 49.658 ;
      RECT 68.63 49.527 69.476 49.612 ;
      RECT 68.676 49.481 69.522 49.566 ;
      RECT 68.722 49.435 69.568 49.52 ;
      RECT 68.768 49.389 69.614 49.474 ;
      RECT 68.814 49.343 69.66 49.428 ;
      RECT 68.86 49.297 69.706 49.382 ;
      RECT 68.906 49.251 69.752 49.336 ;
      RECT 68.952 49.205 69.798 49.29 ;
      RECT 68.998 49.159 69.844 49.244 ;
      RECT 69.044 49.113 69.89 49.198 ;
      RECT 69.09 49.067 69.936 49.152 ;
      RECT 69.136 49.021 69.982 49.106 ;
      RECT 69.182 48.975 70.028 49.06 ;
      RECT 69.228 48.929 70.074 49.014 ;
      RECT 69.274 48.883 70.12 48.968 ;
      RECT 70.102 48.072 70.12 48.968 ;
      RECT 69.32 48.837 70.166 48.922 ;
      RECT 70.115 48.042 70.166 48.922 ;
      RECT 69.366 48.791 70.212 48.876 ;
      RECT 70.161 47.996 70.212 48.876 ;
      RECT 69.412 48.745 70.258 48.83 ;
      RECT 70.207 47.95 70.258 48.83 ;
      RECT 69.458 48.699 70.304 48.784 ;
      RECT 70.253 47.904 70.304 48.784 ;
      RECT 69.504 48.653 70.35 48.738 ;
      RECT 70.299 47.858 70.35 48.738 ;
      RECT 69.55 48.607 70.396 48.692 ;
      RECT 70.345 47.812 70.396 48.692 ;
      RECT 69.596 48.561 70.442 48.646 ;
      RECT 70.391 47.766 70.442 48.646 ;
      RECT 69.642 48.515 70.488 48.6 ;
      RECT 70.437 47.72 70.488 48.6 ;
      RECT 69.688 48.469 70.534 48.554 ;
      RECT 70.483 47.674 70.534 48.554 ;
      RECT 69.734 48.423 70.58 48.508 ;
      RECT 70.529 47.628 70.58 48.508 ;
      RECT 69.78 48.377 70.626 48.462 ;
      RECT 70.575 47.582 70.626 48.462 ;
      RECT 69.826 48.331 70.672 48.416 ;
      RECT 70.621 47.536 70.672 48.416 ;
      RECT 69.872 48.285 70.718 48.37 ;
      RECT 70.667 47.49 70.718 48.37 ;
      RECT 69.918 48.239 70.764 48.324 ;
      RECT 70.713 47.444 70.764 48.324 ;
      RECT 69.964 48.193 70.81 48.278 ;
      RECT 70.759 47.398 70.81 48.278 ;
      RECT 70.01 48.147 70.856 48.232 ;
      RECT 70.805 47.352 70.856 48.232 ;
      RECT 70.056 48.101 70.902 48.186 ;
      RECT 70.851 47.306 70.902 48.186 ;
      RECT 70.897 47.26 70.948 48.14 ;
      RECT 70.943 47.214 70.994 48.094 ;
      RECT 70.989 47.168 71.04 48.048 ;
      RECT 71.035 47.122 71.086 48.002 ;
      RECT 71.081 47.076 71.132 47.956 ;
      RECT 71.127 47.03 71.178 47.91 ;
      RECT 71.173 46.984 71.224 47.864 ;
      RECT 71.219 46.938 71.27 47.818 ;
      RECT 71.265 46.892 71.316 47.772 ;
      RECT 71.311 46.846 71.362 47.726 ;
      RECT 71.357 46.8 71.408 47.68 ;
      RECT 71.403 46.754 71.454 47.634 ;
      RECT 71.449 46.708 71.5 47.588 ;
      RECT 71.495 46.662 71.546 47.542 ;
      RECT 71.541 46.616 71.592 47.496 ;
      RECT 71.587 46.57 71.638 47.45 ;
      RECT 71.633 46.524 71.684 47.404 ;
      RECT 71.679 46.478 71.73 47.358 ;
      RECT 71.725 46.432 71.776 47.312 ;
      RECT 71.771 46.386 71.822 47.266 ;
      RECT 71.817 46.34 71.868 47.22 ;
      RECT 71.863 46.294 71.914 47.174 ;
      RECT 71.909 46.248 71.96 47.128 ;
      RECT 71.955 46.202 72.006 47.082 ;
      RECT 72.001 46.156 72.052 47.036 ;
      RECT 72.047 46.11 72.098 46.99 ;
      RECT 72.093 46.064 72.144 46.944 ;
      RECT 72.139 46.018 72.19 46.898 ;
      RECT 72.185 45.972 72.236 46.852 ;
      RECT 72.231 45.926 72.282 46.806 ;
      RECT 72.277 45.88 72.328 46.76 ;
      RECT 72.323 45.834 72.374 46.714 ;
      RECT 72.369 45.788 72.42 46.668 ;
      RECT 72.415 45.742 72.466 46.622 ;
      RECT 72.461 45.696 72.512 46.576 ;
      RECT 72.507 45.65 72.558 46.53 ;
      RECT 72.553 45.604 72.604 46.484 ;
      RECT 72.599 45.558 72.65 46.438 ;
      RECT 72.645 45.512 72.696 46.392 ;
      RECT 72.691 45.466 72.742 46.346 ;
      RECT 72.737 45.42 72.788 46.3 ;
      RECT 72.783 45.374 72.834 46.254 ;
      RECT 72.829 45.328 72.88 46.208 ;
      RECT 72.875 45.282 72.926 46.162 ;
      RECT 72.921 45.236 72.972 46.116 ;
      RECT 72.967 45.19 73.018 46.07 ;
      RECT 73.013 45.144 73.064 46.024 ;
      RECT 73.059 45.098 73.11 45.978 ;
      RECT 73.105 45.052 73.156 45.932 ;
      RECT 73.151 45.006 73.202 45.886 ;
      RECT 73.197 44.96 73.248 45.84 ;
      RECT 73.243 44.914 73.294 45.794 ;
      RECT 73.289 44.868 73.34 45.748 ;
      RECT 73.335 44.822 73.386 45.702 ;
      RECT 73.381 44.776 73.432 45.656 ;
      RECT 73.427 44.73 73.478 45.61 ;
      RECT 73.473 44.684 73.524 45.564 ;
      RECT 73.519 44.638 73.57 45.518 ;
      RECT 73.565 44.592 73.616 45.472 ;
      RECT 73.611 44.546 73.662 45.426 ;
      RECT 73.657 44.5 73.708 45.38 ;
      RECT 73.703 44.454 73.754 45.334 ;
      RECT 73.749 44.408 73.8 45.288 ;
      RECT 73.795 44.362 73.846 45.242 ;
      RECT 73.841 44.316 73.892 45.196 ;
      RECT 73.887 44.27 73.938 45.15 ;
      RECT 73.933 44.224 73.984 45.104 ;
      RECT 73.979 44.178 74.03 45.058 ;
      RECT 74.025 44.132 74.076 45.012 ;
      RECT 74.071 44.086 74.122 44.966 ;
      RECT 74.117 44.04 74.168 44.92 ;
      RECT 74.163 43.994 74.214 44.874 ;
      RECT 74.209 43.948 74.26 44.828 ;
      RECT 74.255 43.902 74.306 44.782 ;
      RECT 74.301 43.856 74.352 44.736 ;
      RECT 74.347 43.81 74.398 44.69 ;
      RECT 74.393 43.764 74.444 44.644 ;
      RECT 74.439 43.718 74.49 44.598 ;
      RECT 74.485 43.672 74.536 44.552 ;
      RECT 74.531 43.626 74.582 44.506 ;
      RECT 74.577 43.58 74.628 44.46 ;
      RECT 74.623 43.534 74.674 44.414 ;
      RECT 74.669 43.488 74.72 44.368 ;
      RECT 74.715 43.442 74.766 44.322 ;
      RECT 74.761 43.396 74.812 44.276 ;
      RECT 74.807 43.35 74.858 44.23 ;
      RECT 74.853 43.304 74.904 44.184 ;
      RECT 74.899 43.258 74.95 44.138 ;
      RECT 74.945 43.212 74.996 44.092 ;
      RECT 74.991 43.166 75.042 44.046 ;
      RECT 75.037 43.122 75.088 44 ;
      RECT 75.08 43.1 75.134 43.954 ;
      RECT 75.08 43.1 75.18 43.908 ;
      RECT 75.08 43.1 75.226 43.862 ;
      RECT 75.08 43.1 75.272 43.816 ;
      RECT 75.08 43.1 75.318 43.77 ;
      RECT 75.08 43.1 75.364 43.724 ;
      RECT 75.08 43.1 75.41 43.678 ;
      RECT 75.08 43.1 75.456 43.632 ;
      RECT 75.08 43.1 75.502 43.586 ;
      RECT 75.08 43.1 75.548 43.54 ;
      RECT 29.6 68.307 30.038 68.8 ;
      RECT 29.6 68.307 30.084 68.754 ;
      RECT 29.6 68.307 30.13 68.708 ;
      RECT 29.6 68.307 30.176 68.662 ;
      RECT 29.6 68.307 30.222 68.616 ;
      RECT 29.6 68.307 30.268 68.57 ;
      RECT 29.6 68.307 30.314 68.524 ;
      RECT 29.6 68.307 30.36 68.478 ;
      RECT 29.6 68.307 30.406 68.432 ;
      RECT 29.6 68.307 30.452 68.386 ;
      RECT 29.646 68.261 30.498 68.34 ;
      RECT 29.692 68.215 30.544 68.294 ;
      RECT 29.738 68.169 30.59 68.248 ;
      RECT 29.784 68.123 30.636 68.202 ;
      RECT 29.83 68.077 30.682 68.156 ;
      RECT 29.876 68.031 30.728 68.11 ;
      RECT 29.922 67.985 30.774 68.064 ;
      RECT 29.968 67.939 30.82 68.018 ;
      RECT 30.014 67.893 30.866 67.972 ;
      RECT 30.06 67.847 30.912 67.926 ;
      RECT 30.106 67.801 30.958 67.88 ;
      RECT 30.152 67.755 31.004 67.834 ;
      RECT 30.198 67.709 31.05 67.788 ;
      RECT 30.244 67.663 31.096 67.742 ;
      RECT 30.29 67.617 31.142 67.696 ;
      RECT 30.336 67.571 31.188 67.65 ;
      RECT 30.382 67.525 31.234 67.604 ;
      RECT 30.428 67.479 31.28 67.558 ;
      RECT 30.474 67.433 31.326 67.512 ;
      RECT 30.52 67.387 31.372 67.466 ;
      RECT 30.566 67.341 31.418 67.42 ;
      RECT 30.612 67.295 31.464 67.374 ;
      RECT 30.658 67.249 31.51 67.328 ;
      RECT 30.704 67.203 31.556 67.282 ;
      RECT 30.75 67.157 31.602 67.236 ;
      RECT 30.796 67.111 31.648 67.19 ;
      RECT 30.842 67.065 31.694 67.144 ;
      RECT 30.888 67.019 31.74 67.098 ;
      RECT 30.934 66.973 31.786 67.052 ;
      RECT 30.98 66.927 31.832 67.006 ;
      RECT 31.026 66.881 31.878 66.96 ;
      RECT 31.072 66.835 31.924 66.914 ;
      RECT 31.118 66.789 31.97 66.868 ;
      RECT 31.164 66.743 32.016 66.822 ;
      RECT 31.21 66.697 32.062 66.776 ;
      RECT 31.256 66.651 32.108 66.73 ;
      RECT 31.302 66.605 32.154 66.684 ;
      RECT 31.348 66.559 32.2 66.638 ;
      RECT 31.394 66.513 32.246 66.592 ;
      RECT 31.44 66.467 32.292 66.546 ;
      RECT 31.486 66.421 32.338 66.5 ;
      RECT 31.532 66.375 32.384 66.454 ;
      RECT 31.578 66.329 32.43 66.408 ;
      RECT 31.624 66.283 32.476 66.362 ;
      RECT 31.67 66.237 32.522 66.316 ;
      RECT 31.716 66.191 32.568 66.27 ;
      RECT 31.762 66.145 32.614 66.224 ;
      RECT 31.808 66.099 32.66 66.178 ;
      RECT 31.854 66.053 32.706 66.132 ;
      RECT 31.9 66.007 32.752 66.086 ;
      RECT 31.946 65.961 32.798 66.04 ;
      RECT 31.992 65.915 32.844 65.994 ;
      RECT 32.038 65.869 32.89 65.948 ;
      RECT 32.084 65.823 32.936 65.902 ;
      RECT 32.13 65.777 32.982 65.856 ;
      RECT 32.176 65.731 33.028 65.81 ;
      RECT 32.222 65.685 33.074 65.764 ;
      RECT 32.268 65.639 33.12 65.718 ;
      RECT 32.314 65.593 33.166 65.672 ;
      RECT 32.36 65.547 33.212 65.626 ;
      RECT 32.406 65.501 33.258 65.58 ;
      RECT 32.452 65.455 33.304 65.534 ;
      RECT 32.498 65.409 33.35 65.488 ;
      RECT 32.544 65.363 33.396 65.442 ;
      RECT 32.59 65.317 33.442 65.396 ;
      RECT 32.636 65.271 33.488 65.35 ;
      RECT 32.682 65.225 33.534 65.304 ;
      RECT 32.728 65.179 33.58 65.258 ;
      RECT 32.774 65.133 33.626 65.212 ;
      RECT 32.82 65.087 33.672 65.166 ;
      RECT 32.866 65.041 33.718 65.12 ;
      RECT 32.912 64.995 33.764 65.074 ;
      RECT 32.958 64.949 33.81 65.028 ;
      RECT 33.004 64.903 33.856 64.982 ;
      RECT 33.05 64.857 33.902 64.936 ;
      RECT 33.096 64.811 33.948 64.89 ;
      RECT 33.142 64.765 33.994 64.844 ;
      RECT 33.188 64.719 34.04 64.798 ;
      RECT 33.234 64.673 34.086 64.752 ;
      RECT 33.28 64.627 34.132 64.706 ;
      RECT 33.326 64.581 34.178 64.66 ;
      RECT 33.372 64.535 34.224 64.614 ;
      RECT 33.418 64.489 34.27 64.568 ;
      RECT 33.464 64.443 34.316 64.522 ;
      RECT 33.51 64.397 34.362 64.476 ;
      RECT 33.556 64.351 34.408 64.43 ;
      RECT 33.602 64.305 34.454 64.384 ;
      RECT 33.648 64.259 34.5 64.338 ;
      RECT 33.694 64.213 34.546 64.292 ;
      RECT 33.74 64.167 34.592 64.246 ;
      RECT 33.786 64.121 34.638 64.2 ;
      RECT 33.832 64.075 34.684 64.154 ;
      RECT 33.878 64.029 34.73 64.108 ;
      RECT 33.924 63.983 34.776 64.062 ;
      RECT 33.97 63.937 34.822 64.016 ;
      RECT 34.016 63.891 34.868 63.97 ;
      RECT 34.062 63.845 34.914 63.924 ;
      RECT 34.108 63.799 34.96 63.878 ;
      RECT 34.154 63.753 35.006 63.832 ;
      RECT 34.2 63.707 35.052 63.786 ;
      RECT 34.246 63.661 35.098 63.74 ;
      RECT 34.292 63.615 35.144 63.694 ;
      RECT 34.338 63.569 35.19 63.648 ;
      RECT 34.384 63.523 35.236 63.602 ;
      RECT 34.43 63.477 35.282 63.556 ;
      RECT 34.476 63.431 35.328 63.51 ;
      RECT 34.522 63.385 35.374 63.464 ;
      RECT 34.568 63.339 35.42 63.418 ;
      RECT 34.614 63.293 35.466 63.372 ;
      RECT 34.66 63.247 35.512 63.326 ;
      RECT 34.706 63.201 35.558 63.28 ;
      RECT 34.752 63.155 35.604 63.234 ;
      RECT 34.798 63.109 35.65 63.188 ;
      RECT 34.844 63.063 35.696 63.142 ;
      RECT 34.89 63.017 35.742 63.096 ;
      RECT 34.936 62.971 35.788 63.05 ;
      RECT 34.982 62.925 35.834 63.004 ;
      RECT 35.028 62.879 35.88 62.958 ;
      RECT 35.074 62.833 35.926 62.912 ;
      RECT 35.12 62.787 35.972 62.866 ;
      RECT 35.166 62.741 36.018 62.82 ;
      RECT 35.212 62.695 36.064 62.774 ;
      RECT 35.258 62.649 36.11 62.728 ;
      RECT 35.304 62.603 36.156 62.682 ;
      RECT 35.35 62.557 36.202 62.636 ;
      RECT 35.396 62.511 36.248 62.59 ;
      RECT 35.442 62.465 36.294 62.544 ;
      RECT 35.488 62.419 36.34 62.498 ;
      RECT 35.534 62.373 36.386 62.452 ;
      RECT 35.58 62.327 36.432 62.406 ;
      RECT 35.626 62.281 36.478 62.36 ;
      RECT 35.672 62.235 36.524 62.314 ;
      RECT 35.718 62.189 36.57 62.268 ;
      RECT 35.764 62.143 36.616 62.222 ;
      RECT 35.81 62.097 36.662 62.176 ;
      RECT 35.856 62.051 36.708 62.13 ;
      RECT 35.902 62.005 36.754 62.084 ;
      RECT 35.948 61.959 36.8 62.038 ;
      RECT 35.994 61.913 36.846 61.992 ;
      RECT 36.04 61.867 36.892 61.946 ;
      RECT 36.086 61.821 36.938 61.9 ;
      RECT 36.132 61.775 36.984 61.854 ;
      RECT 36.178 61.729 37.03 61.808 ;
      RECT 36.224 61.683 37.076 61.762 ;
      RECT 36.27 61.637 37.122 61.716 ;
      RECT 36.316 61.591 37.168 61.67 ;
      RECT 36.362 61.545 37.214 61.624 ;
      RECT 36.408 61.499 37.26 61.578 ;
      RECT 36.454 61.453 37.306 61.532 ;
      RECT 36.5 61.407 37.352 61.486 ;
      RECT 36.546 61.361 37.398 61.44 ;
      RECT 36.592 61.315 37.444 61.394 ;
      RECT 36.638 61.269 37.49 61.348 ;
      RECT 36.684 61.223 37.536 61.302 ;
      RECT 36.73 61.177 37.582 61.256 ;
      RECT 36.776 61.131 37.628 61.21 ;
      RECT 36.822 61.085 37.674 61.164 ;
      RECT 36.868 61.039 37.72 61.118 ;
      RECT 36.914 60.993 37.766 61.072 ;
      RECT 36.96 60.947 37.812 61.026 ;
      RECT 37.006 60.901 37.858 60.98 ;
      RECT 37.052 60.855 37.904 60.934 ;
      RECT 37.098 60.809 37.95 60.888 ;
      RECT 37.144 60.763 37.996 60.842 ;
      RECT 37.19 60.717 38.042 60.796 ;
      RECT 37.236 60.671 38.088 60.75 ;
      RECT 37.282 60.625 38.134 60.704 ;
      RECT 37.328 60.579 38.18 60.658 ;
      RECT 37.374 60.533 38.226 60.612 ;
      RECT 37.42 60.487 38.272 60.566 ;
      RECT 37.466 60.441 38.318 60.52 ;
      RECT 37.512 60.395 38.364 60.474 ;
      RECT 37.558 60.349 38.41 60.428 ;
      RECT 37.604 60.303 38.456 60.382 ;
      RECT 37.65 60.257 38.502 60.336 ;
      RECT 37.696 60.211 38.548 60.29 ;
      RECT 37.742 60.165 38.594 60.244 ;
      RECT 37.788 60.119 38.64 60.198 ;
      RECT 37.834 60.073 38.686 60.152 ;
      RECT 37.88 60.027 38.732 60.106 ;
      RECT 37.926 59.981 38.778 60.06 ;
      RECT 37.972 59.935 38.824 60.014 ;
      RECT 38.018 59.889 38.87 59.968 ;
      RECT 38.064 59.843 38.916 59.922 ;
      RECT 38.11 59.797 38.962 59.876 ;
      RECT 38.156 59.751 39.008 59.83 ;
      RECT 38.202 59.705 39.054 59.784 ;
      RECT 38.248 59.659 39.1 59.738 ;
      RECT 38.294 59.613 39.146 59.692 ;
      RECT 38.34 59.567 39.192 59.646 ;
      RECT 38.386 59.521 39.238 59.6 ;
      RECT 38.432 59.475 39.284 59.554 ;
      RECT 38.478 59.429 39.33 59.508 ;
      RECT 38.524 59.383 39.376 59.462 ;
      RECT 38.57 59.337 39.422 59.416 ;
      RECT 38.616 59.291 39.468 59.37 ;
      RECT 38.662 59.245 39.514 59.324 ;
      RECT 38.708 59.199 39.56 59.278 ;
      RECT 38.754 59.153 39.606 59.232 ;
      RECT 38.8 59.107 39.652 59.186 ;
      RECT 38.846 59.061 39.698 59.14 ;
      RECT 38.892 59.015 39.744 59.094 ;
      RECT 38.938 58.969 39.79 59.048 ;
      RECT 38.984 58.923 39.836 59.002 ;
      RECT 39.03 58.877 39.882 58.956 ;
      RECT 39.076 58.831 39.928 58.91 ;
      RECT 39.122 58.785 39.974 58.864 ;
      RECT 39.168 58.739 40.02 58.818 ;
      RECT 39.214 58.693 40.066 58.772 ;
      RECT 39.26 58.647 40.112 58.726 ;
      RECT 39.306 58.601 40.158 58.68 ;
      RECT 39.352 58.555 40.204 58.634 ;
      RECT 39.398 58.509 40.25 58.588 ;
      RECT 39.444 58.463 40.296 58.542 ;
      RECT 39.49 58.417 40.342 58.496 ;
      RECT 39.536 58.371 40.388 58.45 ;
      RECT 39.582 58.325 40.434 58.404 ;
      RECT 39.628 58.279 40.48 58.358 ;
      RECT 39.674 58.233 40.526 58.312 ;
      RECT 39.72 58.187 40.572 58.266 ;
      RECT 39.766 58.141 40.618 58.22 ;
      RECT 39.812 58.095 40.664 58.174 ;
      RECT 39.858 58.049 40.71 58.128 ;
      RECT 39.904 58.003 40.756 58.082 ;
      RECT 39.95 57.957 40.802 58.036 ;
      RECT 39.996 57.911 40.848 57.99 ;
      RECT 40.042 57.865 40.894 57.944 ;
      RECT 40.088 57.819 40.94 57.898 ;
      RECT 40.134 57.773 40.986 57.852 ;
      RECT 40.18 57.727 41.032 57.806 ;
      RECT 40.226 57.681 41.078 57.76 ;
      RECT 40.272 57.635 41.124 57.714 ;
      RECT 40.318 57.589 41.17 57.668 ;
      RECT 40.364 57.543 41.216 57.622 ;
      RECT 40.41 57.497 41.262 57.576 ;
      RECT 40.456 57.451 41.308 57.53 ;
      RECT 40.502 57.405 41.354 57.484 ;
      RECT 40.548 57.359 41.4 57.438 ;
      RECT 40.594 57.313 41.446 57.392 ;
      RECT 40.64 57.267 41.492 57.346 ;
      RECT 40.686 57.221 41.538 57.3 ;
      RECT 40.732 57.175 41.584 57.254 ;
      RECT 40.778 57.129 41.63 57.208 ;
      RECT 40.824 57.083 41.676 57.162 ;
      RECT 40.87 57.037 41.722 57.116 ;
      RECT 40.916 56.991 41.768 57.07 ;
      RECT 40.962 56.945 41.814 57.024 ;
      RECT 41.008 56.899 41.86 56.978 ;
      RECT 41.054 56.853 41.9 56.935 ;
      RECT 41.1 56.807 41.946 56.892 ;
      RECT 41.146 56.761 41.992 56.846 ;
      RECT 41.192 56.715 42.038 56.8 ;
      RECT 41.238 56.669 42.084 56.754 ;
      RECT 41.284 56.623 42.13 56.708 ;
      RECT 41.33 56.577 42.176 56.662 ;
      RECT 41.376 56.531 42.222 56.616 ;
      RECT 41.422 56.485 42.268 56.57 ;
      RECT 41.468 56.439 42.314 56.524 ;
      RECT 41.514 56.393 42.36 56.478 ;
      RECT 41.56 56.347 42.406 56.432 ;
      RECT 41.606 56.301 42.452 56.386 ;
      RECT 41.652 56.255 42.498 56.34 ;
      RECT 41.698 56.209 42.544 56.294 ;
      RECT 41.744 56.163 42.59 56.248 ;
      RECT 41.79 56.117 42.636 56.202 ;
      RECT 41.836 56.071 42.682 56.156 ;
      RECT 41.882 56.025 42.728 56.11 ;
      RECT 41.928 55.979 42.774 56.064 ;
      RECT 41.974 55.933 42.82 56.018 ;
      RECT 42.02 55.887 42.866 55.972 ;
      RECT 42.066 55.841 42.912 55.926 ;
      RECT 42.112 55.795 42.958 55.88 ;
      RECT 42.158 55.749 43.004 55.834 ;
      RECT 42.204 55.703 43.05 55.788 ;
      RECT 42.25 55.657 43.096 55.742 ;
      RECT 42.296 55.611 43.142 55.696 ;
      RECT 42.342 55.565 43.188 55.65 ;
      RECT 42.388 55.519 43.234 55.604 ;
      RECT 42.434 55.473 43.28 55.558 ;
      RECT 42.48 55.427 43.326 55.512 ;
      RECT 42.526 55.381 43.372 55.466 ;
      RECT 42.572 55.335 43.418 55.42 ;
      RECT 42.618 55.289 43.464 55.374 ;
      RECT 42.664 55.243 43.51 55.328 ;
      RECT 42.71 55.197 43.556 55.282 ;
      RECT 42.756 55.151 43.602 55.236 ;
      RECT 42.802 55.105 43.648 55.19 ;
      RECT 42.848 55.059 43.694 55.144 ;
      RECT 42.894 55.013 43.74 55.098 ;
      RECT 42.94 54.967 43.786 55.052 ;
      RECT 42.986 54.921 43.832 55.006 ;
      RECT 43.032 54.875 43.878 54.96 ;
      RECT 43.078 54.829 43.924 54.914 ;
      RECT 43.124 54.783 43.97 54.868 ;
      RECT 43.17 54.737 44.016 54.822 ;
      RECT 43.216 54.691 44.062 54.776 ;
      RECT 43.262 54.645 44.108 54.73 ;
      RECT 43.308 54.599 44.154 54.684 ;
      RECT 43.354 54.553 44.2 54.638 ;
      RECT 43.4 54.507 44.246 54.592 ;
      RECT 43.446 54.461 44.292 54.546 ;
      RECT 43.492 54.415 44.338 54.5 ;
      RECT 43.538 54.369 44.384 54.454 ;
      RECT 43.584 54.323 44.43 54.408 ;
      RECT 43.63 54.277 44.476 54.362 ;
      RECT 43.676 54.231 44.522 54.316 ;
      RECT 43.722 54.185 44.568 54.27 ;
      RECT 43.768 54.139 44.614 54.224 ;
      RECT 43.814 54.093 44.66 54.178 ;
      RECT 43.86 54.047 44.706 54.132 ;
      RECT 43.906 54.001 44.752 54.086 ;
      RECT 43.952 53.955 44.798 54.04 ;
      RECT 43.998 53.909 44.844 53.994 ;
      RECT 44.044 53.863 44.89 53.948 ;
      RECT 44.09 53.817 44.936 53.902 ;
      RECT 44.136 53.771 44.982 53.856 ;
      RECT 44.182 53.725 45.028 53.81 ;
      RECT 44.228 53.679 45.074 53.764 ;
      RECT 44.274 53.633 45.12 53.718 ;
      RECT 44.32 53.587 45.166 53.672 ;
      RECT 44.366 53.541 45.212 53.626 ;
      RECT 44.412 53.495 45.258 53.58 ;
      RECT 44.458 53.449 45.304 53.534 ;
      RECT 44.504 53.403 45.35 53.488 ;
      RECT 44.55 53.357 45.396 53.442 ;
      RECT 44.596 53.311 45.442 53.396 ;
      RECT 44.642 53.265 45.488 53.35 ;
      RECT 44.688 53.219 45.534 53.304 ;
      RECT 44.734 53.173 45.58 53.258 ;
      RECT 44.78 53.127 45.626 53.212 ;
      RECT 44.826 53.081 45.672 53.166 ;
      RECT 44.872 53.035 45.718 53.12 ;
      RECT 44.918 52.989 45.764 53.074 ;
      RECT 44.964 52.943 45.81 53.028 ;
      RECT 45.01 52.897 45.856 52.982 ;
      RECT 45.056 52.851 45.902 52.936 ;
      RECT 45.102 52.805 45.948 52.89 ;
      RECT 45.148 52.759 45.994 52.844 ;
      RECT 45.194 52.713 46.04 52.798 ;
      RECT 45.24 52.667 46.086 52.752 ;
      RECT 45.286 52.621 46.132 52.706 ;
      RECT 45.332 52.575 46.178 52.66 ;
      RECT 45.378 52.529 46.224 52.614 ;
      RECT 45.424 52.483 46.27 52.568 ;
      RECT 45.47 52.437 46.316 52.522 ;
      RECT 45.516 52.391 46.362 52.476 ;
      RECT 45.562 52.345 46.408 52.43 ;
      RECT 45.608 52.299 46.454 52.384 ;
      RECT 45.654 52.253 46.5 52.338 ;
      RECT 45.7 52.207 46.546 52.292 ;
      RECT 45.746 52.161 46.592 52.246 ;
      RECT 45.792 52.115 46.638 52.2 ;
      RECT 45.838 52.069 46.684 52.154 ;
      RECT 45.884 52.023 46.73 52.108 ;
      RECT 45.93 51.977 46.776 52.062 ;
      RECT 45.976 51.931 46.822 52.016 ;
      RECT 46.022 51.885 46.868 51.97 ;
      RECT 46.068 51.839 46.914 51.924 ;
      RECT 46.114 51.793 46.96 51.878 ;
      RECT 46.16 51.747 47.006 51.832 ;
      RECT 46.206 51.701 47.052 51.786 ;
      RECT 46.252 51.655 47.098 51.74 ;
      RECT 46.298 51.609 47.144 51.694 ;
      RECT 46.344 51.563 47.19 51.648 ;
      RECT 46.39 51.517 47.236 51.602 ;
      RECT 46.436 51.471 47.282 51.556 ;
      RECT 46.482 51.425 47.328 51.51 ;
      RECT 46.528 51.379 47.374 51.464 ;
      RECT 46.574 51.333 47.42 51.418 ;
      RECT 46.62 51.287 47.466 51.372 ;
      RECT 46.666 51.241 47.512 51.326 ;
      RECT 46.712 51.195 47.558 51.28 ;
      RECT 46.758 51.149 47.604 51.234 ;
      RECT 46.804 51.103 47.65 51.188 ;
      RECT 46.85 51.057 47.696 51.142 ;
      RECT 46.896 51.011 47.742 51.096 ;
      RECT 46.942 50.965 47.788 51.05 ;
      RECT 46.988 50.919 47.834 51.004 ;
      RECT 47.034 50.873 47.88 50.958 ;
      RECT 47.08 50.827 47.926 50.912 ;
      RECT 47.126 50.781 47.972 50.866 ;
      RECT 47.172 50.735 48.018 50.82 ;
      RECT 47.218 50.689 48.064 50.774 ;
      RECT 47.264 50.643 48.11 50.728 ;
      RECT 47.31 50.597 48.156 50.682 ;
      RECT 47.356 50.551 48.202 50.636 ;
      RECT 47.402 50.505 48.248 50.59 ;
      RECT 47.448 50.459 48.294 50.544 ;
      RECT 47.494 50.413 48.34 50.498 ;
      RECT 47.54 50.367 48.386 50.452 ;
      RECT 47.586 50.321 48.432 50.406 ;
      RECT 47.632 50.275 48.478 50.36 ;
      RECT 47.678 50.229 48.524 50.314 ;
      RECT 47.724 50.183 48.57 50.268 ;
      RECT 47.77 50.137 48.616 50.222 ;
      RECT 47.816 50.091 48.662 50.176 ;
      RECT 47.862 50.045 48.708 50.13 ;
      RECT 47.908 49.999 48.754 50.084 ;
      RECT 47.954 49.953 48.8 50.038 ;
      RECT 48 49.907 48.846 49.992 ;
      RECT 48.046 49.861 48.892 49.946 ;
      RECT 48.092 49.815 48.938 49.9 ;
      RECT 48.138 49.769 48.984 49.854 ;
      RECT 48.184 49.723 49.03 49.808 ;
      RECT 48.23 49.677 49.076 49.762 ;
      RECT 48.276 49.631 49.122 49.716 ;
      RECT 48.322 49.585 49.168 49.67 ;
      RECT 48.368 49.539 49.214 49.624 ;
      RECT 48.414 49.493 49.26 49.578 ;
      RECT 48.46 49.447 49.306 49.532 ;
      RECT 48.506 49.401 49.352 49.486 ;
      RECT 48.552 49.355 49.398 49.44 ;
      RECT 48.598 49.309 49.444 49.394 ;
      RECT 48.644 49.263 49.49 49.348 ;
      RECT 48.69 49.217 49.536 49.302 ;
      RECT 48.736 49.171 49.582 49.256 ;
      RECT 48.782 49.125 49.628 49.21 ;
      RECT 48.828 49.079 49.674 49.164 ;
      RECT 48.874 49.033 49.72 49.118 ;
      RECT 48.92 48.987 49.766 49.072 ;
      RECT 48.966 48.941 49.812 49.026 ;
      RECT 49.012 48.895 49.858 48.98 ;
      RECT 49.058 48.849 49.904 48.934 ;
      RECT 49.104 48.803 49.95 48.888 ;
      RECT 49.15 48.757 49.996 48.842 ;
      RECT 49.196 48.711 50.042 48.796 ;
      RECT 49.242 48.665 50.088 48.75 ;
      RECT 49.288 48.619 50.134 48.704 ;
      RECT 49.334 48.573 50.18 48.658 ;
      RECT 49.38 48.527 50.226 48.612 ;
      RECT 49.426 48.481 50.272 48.566 ;
      RECT 49.472 48.435 50.318 48.52 ;
      RECT 49.518 48.389 50.364 48.474 ;
      RECT 49.564 48.343 50.41 48.428 ;
      RECT 49.61 48.297 50.456 48.382 ;
      RECT 49.656 48.251 50.502 48.336 ;
      RECT 49.702 48.205 50.548 48.29 ;
      RECT 49.748 48.159 50.594 48.244 ;
      RECT 49.794 48.113 50.64 48.198 ;
      RECT 49.84 48.067 50.686 48.152 ;
      RECT 49.886 48.021 50.732 48.106 ;
      RECT 49.932 47.975 50.778 48.06 ;
      RECT 49.978 47.929 50.824 48.014 ;
      RECT 50.024 47.883 50.87 47.968 ;
      RECT 50.07 47.837 50.916 47.922 ;
      RECT 50.116 47.791 50.962 47.876 ;
      RECT 50.162 47.745 51.008 47.83 ;
      RECT 50.208 47.699 51.054 47.784 ;
      RECT 50.254 47.653 51.1 47.738 ;
      RECT 50.3 47.607 51.146 47.692 ;
      RECT 50.346 47.561 51.192 47.646 ;
      RECT 50.392 47.515 51.238 47.6 ;
      RECT 50.438 47.469 51.284 47.554 ;
      RECT 50.484 47.423 51.33 47.508 ;
      RECT 50.53 47.377 51.376 47.462 ;
      RECT 50.576 47.331 51.422 47.416 ;
      RECT 50.622 47.285 51.468 47.37 ;
      RECT 50.668 47.239 51.514 47.324 ;
      RECT 50.714 47.193 51.56 47.278 ;
      RECT 50.76 47.147 51.606 47.232 ;
      RECT 50.806 47.101 51.652 47.186 ;
      RECT 50.852 47.055 51.698 47.14 ;
      RECT 50.898 47.009 51.744 47.094 ;
      RECT 50.944 46.963 51.79 47.048 ;
      RECT 50.99 46.917 51.836 47.002 ;
      RECT 51.036 46.871 51.882 46.956 ;
      RECT 51.082 46.825 51.928 46.91 ;
      RECT 51.128 46.779 51.974 46.864 ;
      RECT 51.174 46.733 52.02 46.818 ;
      RECT 51.22 46.687 52.066 46.772 ;
      RECT 51.266 46.641 52.112 46.726 ;
      RECT 51.312 46.595 52.158 46.68 ;
      RECT 51.358 46.549 52.204 46.634 ;
      RECT 51.404 46.503 52.25 46.588 ;
      RECT 51.45 46.457 52.296 46.542 ;
      RECT 51.496 46.411 52.342 46.496 ;
      RECT 51.542 46.365 52.388 46.45 ;
      RECT 51.588 46.319 52.434 46.404 ;
      RECT 51.634 46.273 52.48 46.358 ;
      RECT 51.68 46.227 52.526 46.312 ;
      RECT 51.726 46.181 52.572 46.266 ;
      RECT 51.772 46.135 52.618 46.22 ;
      RECT 51.818 46.089 52.664 46.174 ;
      RECT 51.864 46.043 52.71 46.128 ;
      RECT 51.91 45.997 52.756 46.082 ;
      RECT 51.956 45.951 52.802 46.036 ;
      RECT 52.002 45.905 52.848 45.99 ;
      RECT 52.048 45.859 52.894 45.944 ;
      RECT 52.094 45.813 52.94 45.898 ;
      RECT 52.14 45.767 52.986 45.852 ;
      RECT 52.186 45.721 53.032 45.806 ;
      RECT 52.232 45.675 53.078 45.76 ;
      RECT 52.278 45.629 53.124 45.714 ;
      RECT 52.324 45.583 53.17 45.668 ;
      RECT 52.37 45.537 53.216 45.622 ;
      RECT 52.416 45.491 53.262 45.576 ;
      RECT 52.462 45.445 53.308 45.53 ;
      RECT 52.508 45.399 53.354 45.484 ;
      RECT 52.554 45.353 53.4 45.438 ;
      RECT 52.6 45.307 53.446 45.392 ;
      RECT 52.646 45.261 53.492 45.346 ;
      RECT 52.692 45.215 53.538 45.3 ;
      RECT 52.738 45.169 53.584 45.254 ;
      RECT 52.784 45.123 53.63 45.208 ;
      RECT 52.83 45.077 53.676 45.162 ;
      RECT 52.876 45.031 53.722 45.116 ;
      RECT 52.922 44.985 53.768 45.07 ;
      RECT 52.968 44.939 53.814 45.024 ;
      RECT 53.014 44.893 53.86 44.978 ;
      RECT 53.06 44.847 53.906 44.932 ;
      RECT 53.106 44.801 53.952 44.886 ;
      RECT 53.152 44.755 53.998 44.84 ;
      RECT 53.198 44.709 54.044 44.794 ;
      RECT 53.244 44.663 54.09 44.748 ;
      RECT 53.29 44.617 54.136 44.702 ;
      RECT 53.336 44.571 54.182 44.656 ;
      RECT 53.382 44.525 54.228 44.61 ;
      RECT 53.428 44.479 54.274 44.564 ;
      RECT 53.474 44.433 54.32 44.518 ;
      RECT 53.52 44.387 54.366 44.472 ;
      RECT 53.566 44.341 54.412 44.426 ;
      RECT 53.612 44.295 54.458 44.38 ;
      RECT 53.658 44.249 54.504 44.334 ;
      RECT 53.704 44.203 54.55 44.288 ;
      RECT 53.75 44.157 54.596 44.242 ;
      RECT 53.796 44.111 54.642 44.196 ;
      RECT 53.842 44.065 54.688 44.15 ;
      RECT 53.888 44.019 54.734 44.104 ;
      RECT 53.934 43.973 54.78 44.058 ;
      RECT 53.98 43.927 54.826 44.012 ;
      RECT 54.026 43.881 54.872 43.966 ;
      RECT 54.072 43.835 54.918 43.92 ;
      RECT 54.118 43.789 54.964 43.874 ;
      RECT 54.164 43.743 55.01 43.828 ;
      RECT 54.21 43.697 55.056 43.782 ;
      RECT 54.256 43.651 55.102 43.736 ;
      RECT 54.302 43.605 55.148 43.69 ;
      RECT 54.348 43.559 55.194 43.644 ;
      RECT 54.394 43.513 55.24 43.598 ;
      RECT 54.44 43.467 55.286 43.552 ;
      RECT 54.486 43.421 55.332 43.506 ;
      RECT 54.532 43.375 55.378 43.46 ;
      RECT 54.578 43.329 55.424 43.414 ;
      RECT 54.624 43.283 55.47 43.368 ;
      RECT 54.67 43.237 55.516 43.322 ;
      RECT 54.716 43.191 55.562 43.276 ;
      RECT 54.762 43.145 55.608 43.23 ;
      RECT 54.808 43.099 55.654 43.184 ;
      RECT 54.854 43.053 55.7 43.138 ;
      RECT 54.9 43.007 55.746 43.092 ;
      RECT 54.946 42.961 55.792 43.046 ;
      RECT 54.992 42.915 55.838 43 ;
      RECT 55.038 42.869 55.884 42.954 ;
      RECT 55.084 42.823 55.93 42.908 ;
      RECT 55.13 42.777 55.976 42.862 ;
      RECT 55.176 42.731 56.022 42.816 ;
      RECT 55.222 42.685 56.068 42.77 ;
      RECT 55.268 42.639 56.114 42.724 ;
      RECT 55.314 42.593 56.16 42.678 ;
      RECT 55.36 42.547 56.206 42.632 ;
      RECT 55.406 42.501 56.252 42.586 ;
      RECT 55.452 42.455 56.298 42.54 ;
      RECT 55.498 42.409 56.344 42.494 ;
      RECT 55.544 42.363 56.39 42.448 ;
      RECT 55.59 42.317 56.436 42.402 ;
      RECT 55.636 42.271 56.482 42.356 ;
      RECT 55.682 42.225 56.528 42.31 ;
      RECT 55.728 42.179 56.574 42.264 ;
      RECT 55.774 42.133 56.62 42.218 ;
      RECT 55.82 42.087 56.666 42.172 ;
      RECT 55.866 42.041 56.712 42.126 ;
      RECT 55.912 41.995 56.758 42.08 ;
      RECT 55.958 41.949 56.804 42.034 ;
      RECT 56.004 41.903 56.85 41.988 ;
      RECT 56.05 41.857 56.896 41.942 ;
      RECT 56.096 41.811 56.942 41.896 ;
      RECT 56.142 41.765 56.988 41.85 ;
      RECT 56.188 41.719 57.034 41.804 ;
      RECT 56.234 41.673 57.08 41.758 ;
      RECT 56.28 41.627 57.126 41.712 ;
      RECT 56.326 41.581 57.172 41.666 ;
      RECT 56.372 41.535 57.218 41.62 ;
      RECT 56.418 41.489 57.264 41.574 ;
      RECT 56.464 41.443 57.31 41.528 ;
      RECT 56.51 41.397 57.356 41.482 ;
      RECT 56.556 41.351 57.402 41.436 ;
      RECT 56.602 41.305 57.448 41.39 ;
      RECT 56.648 41.259 57.494 41.344 ;
      RECT 56.694 41.213 57.54 41.298 ;
      RECT 56.74 41.167 57.586 41.252 ;
      RECT 56.786 41.121 57.632 41.206 ;
      RECT 56.832 41.075 57.678 41.16 ;
      RECT 56.878 41.029 57.724 41.114 ;
      RECT 56.924 40.983 57.77 41.068 ;
      RECT 56.97 40.937 57.816 41.022 ;
      RECT 57.016 40.891 57.862 40.976 ;
      RECT 57.062 40.845 57.908 40.93 ;
      RECT 57.108 40.799 57.954 40.884 ;
      RECT 57.154 40.753 58 40.838 ;
      RECT 57.2 40.707 58.046 40.792 ;
      RECT 57.246 40.661 58.092 40.746 ;
      RECT 57.292 40.615 58.138 40.7 ;
      RECT 57.338 40.569 58.184 40.654 ;
      RECT 57.384 40.523 58.23 40.608 ;
      RECT 57.43 40.477 58.276 40.562 ;
      RECT 57.476 40.431 58.322 40.516 ;
      RECT 57.522 40.385 58.368 40.47 ;
      RECT 57.568 40.339 58.414 40.424 ;
      RECT 57.614 40.293 58.46 40.378 ;
      RECT 57.66 40.247 58.506 40.332 ;
      RECT 57.706 40.201 58.552 40.286 ;
      RECT 57.752 40.155 58.598 40.24 ;
      RECT 57.798 40.109 58.644 40.194 ;
      RECT 57.844 40.063 58.69 40.148 ;
      RECT 57.89 40.017 58.736 40.102 ;
      RECT 57.936 39.971 58.782 40.056 ;
      RECT 57.982 39.925 58.828 40.01 ;
      RECT 58.028 39.879 58.874 39.964 ;
      RECT 58.074 39.833 58.92 39.918 ;
      RECT 58.12 39.787 58.966 39.872 ;
      RECT 58.166 39.741 59.012 39.826 ;
      RECT 58.212 39.695 59.058 39.78 ;
      RECT 58.258 39.649 59.104 39.734 ;
      RECT 58.304 39.603 59.15 39.688 ;
      RECT 58.35 39.557 59.196 39.642 ;
      RECT 58.396 39.511 59.242 39.596 ;
      RECT 58.442 39.465 59.288 39.55 ;
      RECT 58.488 39.419 59.334 39.504 ;
      RECT 58.534 39.373 59.38 39.458 ;
      RECT 58.58 39.327 59.426 39.412 ;
      RECT 58.626 39.281 59.472 39.366 ;
      RECT 58.672 39.235 59.518 39.32 ;
      RECT 58.718 39.189 59.564 39.274 ;
      RECT 58.764 39.143 59.61 39.228 ;
      RECT 58.81 39.097 59.656 39.182 ;
      RECT 58.856 39.051 59.702 39.136 ;
      RECT 58.902 39.005 59.748 39.09 ;
      RECT 58.948 38.959 59.794 39.044 ;
      RECT 58.994 38.913 59.84 38.998 ;
      RECT 59.04 38.867 59.886 38.952 ;
      RECT 59.086 38.821 59.932 38.906 ;
      RECT 59.132 38.775 59.978 38.86 ;
      RECT 59.178 38.729 60.024 38.814 ;
      RECT 59.224 38.683 60.07 38.768 ;
      RECT 59.27 38.637 60.116 38.722 ;
      RECT 59.316 38.591 60.162 38.676 ;
      RECT 59.362 38.545 60.208 38.63 ;
      RECT 59.408 38.499 60.254 38.584 ;
      RECT 59.454 38.453 60.3 38.538 ;
      RECT 59.5 38.407 60.346 38.492 ;
      RECT 59.546 38.361 60.392 38.446 ;
      RECT 59.592 38.315 60.438 38.4 ;
      RECT 59.638 38.269 60.484 38.354 ;
      RECT 59.684 38.223 60.53 38.308 ;
      RECT 59.73 38.177 60.576 38.262 ;
      RECT 59.776 38.131 60.622 38.216 ;
      RECT 59.822 38.085 60.668 38.17 ;
      RECT 59.868 38.039 60.714 38.124 ;
      RECT 59.914 37.993 60.76 38.078 ;
      RECT 59.96 37.947 60.806 38.032 ;
      RECT 60.006 37.901 60.852 37.986 ;
      RECT 60.052 37.855 60.898 37.94 ;
      RECT 60.098 37.809 60.944 37.894 ;
      RECT 60.144 37.763 60.99 37.848 ;
      RECT 60.19 37.717 61.036 37.802 ;
      RECT 60.236 37.671 61.082 37.756 ;
      RECT 60.282 37.625 61.128 37.71 ;
      RECT 60.328 37.579 61.174 37.664 ;
      RECT 60.374 37.533 61.22 37.618 ;
      RECT 60.42 37.487 61.266 37.572 ;
      RECT 60.466 37.441 61.312 37.526 ;
      RECT 60.512 37.395 61.358 37.48 ;
      RECT 60.558 37.349 61.404 37.434 ;
      RECT 60.604 37.303 61.45 37.388 ;
      RECT 60.65 37.257 61.496 37.342 ;
      RECT 60.696 37.211 61.542 37.296 ;
      RECT 60.742 37.165 61.588 37.25 ;
      RECT 60.788 37.119 61.634 37.204 ;
      RECT 60.834 37.073 61.68 37.158 ;
      RECT 60.88 37.027 61.726 37.112 ;
      RECT 60.926 36.981 61.772 37.066 ;
      RECT 60.972 36.935 61.818 37.02 ;
      RECT 61.018 36.889 61.864 36.974 ;
      RECT 61.064 36.843 61.91 36.928 ;
      RECT 61.11 36.797 61.956 36.882 ;
      RECT 61.156 36.751 62.002 36.836 ;
      RECT 61.202 36.705 62.048 36.79 ;
      RECT 61.248 36.659 62.094 36.744 ;
      RECT 61.294 36.613 62.14 36.698 ;
      RECT 61.34 36.567 62.186 36.652 ;
      RECT 61.386 36.521 62.232 36.606 ;
      RECT 61.432 36.475 62.278 36.56 ;
      RECT 61.478 36.429 62.324 36.514 ;
      RECT 61.524 36.383 62.37 36.468 ;
      RECT 61.57 36.337 62.416 36.422 ;
      RECT 61.616 36.291 62.462 36.376 ;
      RECT 61.662 36.245 62.508 36.33 ;
      RECT 61.708 36.199 62.554 36.284 ;
      RECT 61.754 36.153 62.6 36.238 ;
      RECT 61.8 36.107 62.646 36.192 ;
      RECT 61.846 36.061 62.692 36.146 ;
      RECT 61.892 36.015 62.738 36.1 ;
      RECT 61.938 35.969 62.784 36.054 ;
      RECT 61.984 35.923 62.83 36.008 ;
      RECT 62.03 35.877 62.876 35.962 ;
      RECT 62.076 35.831 62.922 35.916 ;
      RECT 62.122 35.785 62.968 35.87 ;
      RECT 62.168 35.739 63.014 35.824 ;
      RECT 62.214 35.693 63.06 35.778 ;
      RECT 62.26 35.647 63.106 35.732 ;
      RECT 62.306 35.601 63.152 35.686 ;
      RECT 62.352 35.555 63.198 35.64 ;
      RECT 62.398 35.509 63.244 35.594 ;
      RECT 62.444 35.463 63.29 35.548 ;
      RECT 62.49 35.417 63.336 35.502 ;
      RECT 62.536 35.371 63.382 35.456 ;
      RECT 63.364 34.566 63.382 35.456 ;
      RECT 62.582 35.325 63.428 35.41 ;
      RECT 63.365 34.542 63.428 35.41 ;
      RECT 62.628 35.279 63.474 35.364 ;
      RECT 63.411 34.496 63.474 35.364 ;
      RECT 62.674 35.233 63.52 35.318 ;
      RECT 63.457 34.45 63.52 35.318 ;
      RECT 62.72 35.187 63.566 35.272 ;
      RECT 63.503 34.404 63.566 35.272 ;
      RECT 62.766 35.141 63.612 35.226 ;
      RECT 63.549 34.358 63.612 35.226 ;
      RECT 62.812 35.095 63.658 35.18 ;
      RECT 63.595 34.312 63.658 35.18 ;
      RECT 62.858 35.049 63.704 35.134 ;
      RECT 63.641 34.266 63.704 35.134 ;
      RECT 62.904 35.003 63.75 35.088 ;
      RECT 63.687 34.22 63.75 35.088 ;
      RECT 62.95 34.957 63.796 35.042 ;
      RECT 63.733 34.174 63.796 35.042 ;
      RECT 62.996 34.911 63.842 34.996 ;
      RECT 63.779 34.128 63.842 34.996 ;
      RECT 63.042 34.865 63.888 34.95 ;
      RECT 63.825 34.082 63.888 34.95 ;
      RECT 63.088 34.819 63.934 34.904 ;
      RECT 63.871 34.036 63.934 34.904 ;
      RECT 63.134 34.773 63.98 34.858 ;
      RECT 63.917 33.99 63.98 34.858 ;
      RECT 63.18 34.727 64.026 34.812 ;
      RECT 63.963 33.944 64.026 34.812 ;
      RECT 63.226 34.681 64.072 34.766 ;
      RECT 64.009 33.898 64.072 34.766 ;
      RECT 63.272 34.635 64.118 34.72 ;
      RECT 64.055 33.852 64.118 34.72 ;
      RECT 63.318 34.589 64.164 34.674 ;
      RECT 64.101 33.806 64.164 34.674 ;
      RECT 64.147 33.76 64.21 34.628 ;
      RECT 64.193 33.714 64.256 34.582 ;
      RECT 64.239 33.668 64.302 34.536 ;
      RECT 64.285 33.622 64.348 34.49 ;
      RECT 64.331 33.576 64.394 34.444 ;
      RECT 64.377 33.53 64.44 34.398 ;
      RECT 64.423 33.484 64.486 34.352 ;
      RECT 64.469 33.438 64.532 34.306 ;
      RECT 64.515 33.392 64.578 34.26 ;
      RECT 64.561 33.346 64.624 34.214 ;
      RECT 64.607 33.3 64.67 34.168 ;
      RECT 64.653 33.254 64.716 34.122 ;
      RECT 64.699 33.208 64.762 34.076 ;
      RECT 64.745 33.162 64.808 34.03 ;
      RECT 64.791 33.116 64.854 33.984 ;
      RECT 64.837 33.07 64.9 33.938 ;
      RECT 64.883 33.024 64.946 33.892 ;
      RECT 64.929 32.978 64.992 33.846 ;
      RECT 64.975 32.932 65.038 33.8 ;
      RECT 65.021 32.886 65.084 33.754 ;
      RECT 65.067 32.84 65.13 33.708 ;
      RECT 65.113 32.794 65.176 33.662 ;
      RECT 65.159 32.748 65.222 33.616 ;
      RECT 65.205 32.702 65.268 33.57 ;
      RECT 65.251 32.656 65.314 33.524 ;
      RECT 65.297 32.61 65.36 33.478 ;
      RECT 65.343 32.564 65.406 33.432 ;
      RECT 65.389 32.518 65.452 33.386 ;
      RECT 65.435 32.472 65.498 33.34 ;
      RECT 65.481 32.426 65.544 33.294 ;
      RECT 65.527 32.38 65.59 33.248 ;
      RECT 65.573 32.334 65.636 33.202 ;
      RECT 65.619 32.288 65.682 33.156 ;
      RECT 65.665 32.242 65.728 33.11 ;
      RECT 65.711 32.196 65.774 33.064 ;
      RECT 65.757 32.15 65.82 33.018 ;
      RECT 65.803 32.104 65.866 32.972 ;
      RECT 65.849 32.058 65.912 32.926 ;
      RECT 65.895 32.012 65.958 32.88 ;
      RECT 65.941 31.966 66.004 32.834 ;
      RECT 65.987 31.92 66.05 32.788 ;
      RECT 66.033 31.874 66.096 32.742 ;
      RECT 66.079 31.828 66.142 32.696 ;
      RECT 66.125 31.782 66.188 32.65 ;
      RECT 66.171 31.736 66.234 32.604 ;
      RECT 66.217 31.69 66.28 32.558 ;
      RECT 66.263 31.644 66.326 32.512 ;
      RECT 66.309 31.598 66.372 32.466 ;
      RECT 66.355 31.552 66.418 32.42 ;
      RECT 66.401 31.506 66.464 32.374 ;
      RECT 66.447 31.46 66.51 32.328 ;
      RECT 66.493 31.414 66.556 32.282 ;
      RECT 66.539 31.368 66.602 32.236 ;
      RECT 66.585 31.322 66.648 32.19 ;
      RECT 66.631 31.276 66.694 32.144 ;
      RECT 66.677 31.23 66.74 32.098 ;
      RECT 66.723 31.184 66.786 32.052 ;
      RECT 66.769 31.138 66.832 32.006 ;
      RECT 66.815 31.092 66.878 31.96 ;
      RECT 66.861 31.046 66.924 31.914 ;
      RECT 66.907 31 66.97 31.868 ;
      RECT 66.953 30.954 67.016 31.822 ;
      RECT 66.999 30.908 67.062 31.776 ;
      RECT 67.045 30.862 67.108 31.73 ;
      RECT 67.091 30.816 67.154 31.684 ;
      RECT 67.137 30.77 67.2 31.638 ;
      RECT 67.183 30.724 67.246 31.592 ;
      RECT 67.229 30.678 67.292 31.546 ;
      RECT 67.275 30.632 67.338 31.5 ;
      RECT 67.321 30.586 67.384 31.454 ;
      RECT 67.367 30.54 67.43 31.408 ;
      RECT 67.413 30.494 67.476 31.362 ;
      RECT 67.459 30.448 67.522 31.316 ;
      RECT 67.505 30.402 67.568 31.27 ;
      RECT 67.551 30.356 67.614 31.224 ;
      RECT 67.597 30.31 67.66 31.178 ;
      RECT 67.643 30.264 67.706 31.132 ;
      RECT 67.689 30.218 67.752 31.086 ;
      RECT 67.735 30.172 67.798 31.04 ;
      RECT 67.781 30.126 67.844 30.994 ;
      RECT 67.827 30.08 67.89 30.948 ;
      RECT 67.873 30.034 67.936 30.902 ;
      RECT 67.919 29.988 67.982 30.856 ;
      RECT 67.965 29.942 68.028 30.81 ;
      RECT 68.011 29.896 68.074 30.764 ;
      RECT 68.057 29.85 68.12 30.718 ;
      RECT 68.103 29.804 68.166 30.672 ;
      RECT 68.149 29.758 68.212 30.626 ;
      RECT 68.195 29.712 68.258 30.58 ;
      RECT 68.241 29.666 68.304 30.534 ;
      RECT 68.287 29.622 68.35 30.488 ;
      RECT 68.33 29.6 68.396 30.442 ;
      RECT 68.33 29.6 68.442 30.396 ;
      RECT 68.33 29.6 68.488 30.35 ;
      RECT 68.33 29.6 68.534 30.304 ;
      RECT 68.33 29.6 68.58 30.258 ;
      RECT 68.33 29.6 68.626 30.212 ;
      RECT 68.33 29.6 68.672 30.166 ;
      RECT 68.33 29.6 68.718 30.12 ;
      RECT 68.33 29.6 68.764 30.074 ;
      RECT 68.33 29.6 68.81 30.028 ;
      RECT 16.1 61.557 16.538 62.05 ;
      RECT 16.1 61.557 16.584 62.004 ;
      RECT 16.1 61.557 16.63 61.958 ;
      RECT 16.1 61.557 16.676 61.912 ;
      RECT 16.1 61.557 16.722 61.866 ;
      RECT 16.1 61.557 16.768 61.82 ;
      RECT 16.1 61.557 16.814 61.774 ;
      RECT 16.1 61.557 16.86 61.728 ;
      RECT 16.1 61.557 16.906 61.682 ;
      RECT 16.1 61.557 16.952 61.636 ;
      RECT 16.146 61.511 16.998 61.59 ;
      RECT 16.928 60.729 16.998 61.59 ;
      RECT 16.192 61.465 17.044 61.544 ;
      RECT 16.974 60.683 17.044 61.544 ;
      RECT 16.238 61.419 17.09 61.498 ;
      RECT 17.02 60.637 17.09 61.498 ;
      RECT 16.284 61.373 17.136 61.452 ;
      RECT 17.066 60.591 17.136 61.452 ;
      RECT 16.33 61.327 17.182 61.406 ;
      RECT 17.112 60.545 17.182 61.406 ;
      RECT 16.376 61.281 17.228 61.36 ;
      RECT 17.158 60.499 17.228 61.36 ;
      RECT 16.422 61.235 17.274 61.314 ;
      RECT 17.204 60.453 17.274 61.314 ;
      RECT 16.468 61.189 17.32 61.268 ;
      RECT 17.25 60.407 17.32 61.268 ;
      RECT 16.514 61.143 17.366 61.222 ;
      RECT 17.296 60.361 17.366 61.222 ;
      RECT 16.56 61.097 17.412 61.176 ;
      RECT 17.342 60.315 17.412 61.176 ;
      RECT 16.606 61.051 17.458 61.13 ;
      RECT 17.388 60.269 17.458 61.13 ;
      RECT 16.652 61.005 17.504 61.084 ;
      RECT 17.434 60.223 17.504 61.084 ;
      RECT 16.698 60.959 17.55 61.038 ;
      RECT 17.48 60.177 17.55 61.038 ;
      RECT 16.744 60.913 17.596 60.992 ;
      RECT 17.526 60.131 17.596 60.992 ;
      RECT 16.79 60.867 17.642 60.946 ;
      RECT 17.572 60.085 17.642 60.946 ;
      RECT 16.836 60.821 17.688 60.9 ;
      RECT 17.618 60.039 17.688 60.9 ;
      RECT 16.882 60.775 17.734 60.854 ;
      RECT 17.664 59.993 17.734 60.854 ;
      RECT 17.71 59.947 17.78 60.808 ;
      RECT 17.756 59.901 17.826 60.762 ;
      RECT 17.802 59.855 17.872 60.716 ;
      RECT 17.848 59.809 17.918 60.67 ;
      RECT 17.894 59.763 17.964 60.624 ;
      RECT 17.94 59.717 18.01 60.578 ;
      RECT 17.986 59.671 18.056 60.532 ;
      RECT 18.032 59.625 18.102 60.486 ;
      RECT 18.078 59.579 18.148 60.44 ;
      RECT 18.124 59.533 18.194 60.394 ;
      RECT 18.17 59.487 18.24 60.348 ;
      RECT 18.216 59.441 18.286 60.302 ;
      RECT 18.262 59.395 18.332 60.256 ;
      RECT 18.308 59.349 18.378 60.21 ;
      RECT 18.354 59.303 18.424 60.164 ;
      RECT 18.4 59.257 18.47 60.118 ;
      RECT 18.446 59.211 18.516 60.072 ;
      RECT 18.492 59.165 18.562 60.026 ;
      RECT 18.538 59.119 18.608 59.98 ;
      RECT 18.584 59.073 18.654 59.934 ;
      RECT 18.63 59.027 18.7 59.888 ;
      RECT 18.676 58.981 18.746 59.842 ;
      RECT 18.722 58.935 18.792 59.796 ;
      RECT 18.768 58.889 18.838 59.75 ;
      RECT 18.814 58.843 18.884 59.704 ;
      RECT 18.86 58.797 18.93 59.658 ;
      RECT 18.906 58.751 18.976 59.612 ;
      RECT 18.952 58.705 19.022 59.566 ;
      RECT 18.998 58.659 19.068 59.52 ;
      RECT 19.044 58.613 19.114 59.474 ;
      RECT 19.09 58.567 19.16 59.428 ;
      RECT 19.136 58.521 19.206 59.382 ;
      RECT 19.182 58.475 19.252 59.336 ;
      RECT 19.228 58.429 19.298 59.29 ;
      RECT 19.274 58.383 19.344 59.244 ;
      RECT 19.32 58.337 19.39 59.198 ;
      RECT 19.366 58.291 19.436 59.152 ;
      RECT 19.412 58.245 19.482 59.106 ;
      RECT 19.458 58.199 19.528 59.06 ;
      RECT 19.504 58.153 19.574 59.014 ;
      RECT 19.55 58.107 19.62 58.968 ;
      RECT 19.596 58.061 19.666 58.922 ;
      RECT 19.642 58.015 19.712 58.876 ;
      RECT 19.688 57.969 19.758 58.83 ;
      RECT 19.734 57.923 19.804 58.784 ;
      RECT 19.78 57.877 19.85 58.738 ;
      RECT 19.826 57.831 19.896 58.692 ;
      RECT 19.872 57.785 19.942 58.646 ;
      RECT 19.918 57.739 19.988 58.6 ;
      RECT 19.964 57.693 20.034 58.554 ;
      RECT 20.01 57.647 20.08 58.508 ;
      RECT 20.056 57.601 20.126 58.462 ;
      RECT 20.102 57.555 20.172 58.416 ;
      RECT 20.148 57.509 20.218 58.37 ;
      RECT 20.194 57.463 20.264 58.324 ;
      RECT 20.24 57.417 20.31 58.278 ;
      RECT 20.286 57.371 20.356 58.232 ;
      RECT 20.332 57.325 20.402 58.186 ;
      RECT 20.378 57.279 20.448 58.14 ;
      RECT 20.424 57.233 20.494 58.094 ;
      RECT 20.47 57.187 20.54 58.048 ;
      RECT 20.516 57.141 20.586 58.002 ;
      RECT 20.562 57.095 20.632 57.956 ;
      RECT 20.608 57.049 20.678 57.91 ;
      RECT 20.654 57.003 20.724 57.864 ;
      RECT 20.7 56.957 20.77 57.818 ;
      RECT 20.746 56.911 20.816 57.772 ;
      RECT 20.792 56.865 20.862 57.726 ;
      RECT 20.838 56.819 20.908 57.68 ;
      RECT 20.884 56.773 20.954 57.634 ;
      RECT 20.93 56.727 21 57.588 ;
      RECT 20.976 56.681 21.046 57.542 ;
      RECT 21.022 56.635 21.092 57.496 ;
      RECT 21.068 56.589 21.138 57.45 ;
      RECT 21.114 56.543 21.184 57.404 ;
      RECT 21.16 56.497 21.23 57.358 ;
      RECT 21.206 56.451 21.276 57.312 ;
      RECT 21.252 56.405 21.322 57.266 ;
      RECT 21.298 56.359 21.368 57.22 ;
      RECT 21.344 56.313 21.414 57.174 ;
      RECT 21.39 56.267 21.46 57.128 ;
      RECT 21.436 56.221 21.506 57.082 ;
      RECT 21.482 56.175 21.552 57.036 ;
      RECT 21.528 56.129 21.598 56.99 ;
      RECT 21.574 56.083 21.644 56.944 ;
      RECT 21.62 56.037 21.69 56.898 ;
      RECT 21.666 55.991 21.736 56.852 ;
      RECT 21.712 55.945 21.782 56.806 ;
      RECT 21.758 55.899 21.828 56.76 ;
      RECT 21.804 55.853 21.874 56.714 ;
      RECT 21.85 55.807 21.92 56.668 ;
      RECT 21.896 55.761 21.966 56.622 ;
      RECT 21.942 55.715 22.012 56.576 ;
      RECT 21.988 55.669 22.058 56.53 ;
      RECT 22.034 55.623 22.104 56.484 ;
      RECT 22.08 55.577 22.15 56.438 ;
      RECT 22.126 55.531 22.196 56.392 ;
      RECT 22.172 55.485 22.242 56.346 ;
      RECT 22.218 55.439 22.288 56.3 ;
      RECT 22.264 55.393 22.334 56.254 ;
      RECT 22.31 55.347 22.38 56.208 ;
      RECT 22.356 55.301 22.426 56.162 ;
      RECT 22.402 55.255 22.472 56.116 ;
      RECT 22.448 55.209 22.518 56.07 ;
      RECT 22.494 55.163 22.564 56.024 ;
      RECT 22.54 55.117 22.61 55.978 ;
      RECT 22.586 55.071 22.656 55.932 ;
      RECT 22.632 55.025 22.702 55.886 ;
      RECT 22.678 54.979 22.748 55.84 ;
      RECT 22.724 54.933 22.794 55.794 ;
      RECT 22.77 54.887 22.84 55.748 ;
      RECT 22.816 54.841 22.886 55.702 ;
      RECT 22.862 54.795 22.932 55.656 ;
      RECT 22.908 54.749 22.978 55.61 ;
      RECT 22.954 54.703 23.024 55.564 ;
      RECT 23 54.657 23.07 55.518 ;
      RECT 23.046 54.611 23.116 55.472 ;
      RECT 23.092 54.565 23.162 55.426 ;
      RECT 23.138 54.519 23.208 55.38 ;
      RECT 23.184 54.473 23.254 55.334 ;
      RECT 23.23 54.427 23.3 55.288 ;
      RECT 23.276 54.381 23.346 55.242 ;
      RECT 23.322 54.335 23.392 55.196 ;
      RECT 23.368 54.289 23.438 55.15 ;
      RECT 23.414 54.243 23.484 55.104 ;
      RECT 23.46 54.197 23.53 55.058 ;
      RECT 23.506 54.151 23.576 55.012 ;
      RECT 23.552 54.105 23.622 54.966 ;
      RECT 23.598 54.059 23.668 54.92 ;
      RECT 23.644 54.013 23.714 54.874 ;
      RECT 23.69 53.967 23.76 54.828 ;
      RECT 23.736 53.921 23.806 54.782 ;
      RECT 23.782 53.875 23.852 54.736 ;
      RECT 23.828 53.829 23.898 54.69 ;
      RECT 23.874 53.783 23.944 54.644 ;
      RECT 23.92 53.737 23.99 54.598 ;
      RECT 23.966 53.691 24.036 54.552 ;
      RECT 24.012 53.645 24.082 54.506 ;
      RECT 24.058 53.599 24.128 54.46 ;
      RECT 24.104 53.553 24.174 54.414 ;
      RECT 24.15 53.507 24.22 54.368 ;
      RECT 24.196 53.461 24.266 54.322 ;
      RECT 24.242 53.415 24.312 54.276 ;
      RECT 24.288 53.369 24.358 54.23 ;
      RECT 24.334 53.323 24.404 54.184 ;
      RECT 24.38 53.277 24.45 54.138 ;
      RECT 24.426 53.231 24.496 54.092 ;
      RECT 24.472 53.185 24.542 54.046 ;
      RECT 24.518 53.139 24.588 54 ;
      RECT 24.564 53.093 24.634 53.954 ;
      RECT 24.61 53.047 24.68 53.908 ;
      RECT 24.656 53.001 24.726 53.862 ;
      RECT 24.702 52.955 24.772 53.816 ;
      RECT 24.748 52.909 24.818 53.77 ;
      RECT 24.794 52.863 24.864 53.724 ;
      RECT 24.84 52.817 24.91 53.678 ;
      RECT 24.886 52.771 24.956 53.632 ;
      RECT 24.932 52.725 25.002 53.586 ;
      RECT 24.978 52.679 25.048 53.54 ;
      RECT 25.024 52.633 25.094 53.494 ;
      RECT 25.07 52.587 25.14 53.448 ;
      RECT 25.116 52.541 25.186 53.402 ;
      RECT 25.162 52.495 25.232 53.356 ;
      RECT 25.208 52.449 25.278 53.31 ;
      RECT 25.254 52.403 25.324 53.264 ;
      RECT 25.3 52.357 25.37 53.218 ;
      RECT 25.346 52.311 25.416 53.172 ;
      RECT 25.392 52.265 25.462 53.126 ;
      RECT 25.438 52.219 25.508 53.08 ;
      RECT 25.484 52.173 25.554 53.034 ;
      RECT 25.53 52.127 25.6 52.988 ;
      RECT 25.576 52.081 25.646 52.942 ;
      RECT 25.622 52.035 25.692 52.896 ;
      RECT 25.668 51.989 25.738 52.85 ;
      RECT 25.714 51.943 25.784 52.804 ;
      RECT 25.76 51.897 25.83 52.758 ;
      RECT 25.806 51.851 25.876 52.712 ;
      RECT 25.852 51.805 25.922 52.666 ;
      RECT 25.898 51.759 25.968 52.62 ;
      RECT 25.944 51.713 26.014 52.574 ;
      RECT 25.99 51.667 26.06 52.528 ;
      RECT 26.036 51.621 26.106 52.482 ;
      RECT 26.082 51.575 26.152 52.436 ;
      RECT 26.128 51.529 26.198 52.39 ;
      RECT 26.174 51.483 26.244 52.344 ;
      RECT 26.22 51.437 26.29 52.298 ;
      RECT 26.266 51.391 26.336 52.252 ;
      RECT 26.312 51.345 26.382 52.206 ;
      RECT 26.358 51.299 26.428 52.16 ;
      RECT 26.404 51.253 26.474 52.114 ;
      RECT 26.45 51.207 26.52 52.068 ;
      RECT 26.496 51.161 26.566 52.022 ;
      RECT 26.542 51.115 26.612 51.976 ;
      RECT 26.588 51.069 26.658 51.93 ;
      RECT 26.634 51.023 26.704 51.884 ;
      RECT 26.68 50.977 26.75 51.838 ;
      RECT 26.726 50.931 26.796 51.792 ;
      RECT 26.772 50.885 26.842 51.746 ;
      RECT 26.818 50.839 26.888 51.7 ;
      RECT 26.864 50.793 26.934 51.654 ;
      RECT 26.91 50.747 26.98 51.608 ;
      RECT 26.956 50.701 27.026 51.562 ;
      RECT 27.002 50.655 27.072 51.516 ;
      RECT 27.048 50.609 27.118 51.47 ;
      RECT 27.094 50.563 27.164 51.424 ;
      RECT 27.14 50.517 27.21 51.378 ;
      RECT 27.186 50.471 27.256 51.332 ;
      RECT 27.232 50.425 27.302 51.286 ;
      RECT 27.278 50.379 27.348 51.24 ;
      RECT 27.324 50.333 27.394 51.194 ;
      RECT 27.37 50.287 27.44 51.148 ;
      RECT 27.416 50.241 27.486 51.102 ;
      RECT 27.462 50.195 27.532 51.056 ;
      RECT 27.508 50.149 27.578 51.01 ;
      RECT 27.554 50.103 27.624 50.964 ;
      RECT 27.6 50.057 27.67 50.918 ;
      RECT 27.646 50.011 27.716 50.872 ;
      RECT 27.692 49.965 27.762 50.826 ;
      RECT 27.738 49.919 27.808 50.78 ;
      RECT 27.784 49.873 27.854 50.734 ;
      RECT 27.83 49.827 27.9 50.688 ;
      RECT 27.876 49.781 27.946 50.642 ;
      RECT 27.922 49.735 27.992 50.596 ;
      RECT 27.968 49.689 28.038 50.55 ;
      RECT 28.014 49.643 28.084 50.504 ;
      RECT 28.06 49.597 28.13 50.458 ;
      RECT 28.106 49.551 28.176 50.412 ;
      RECT 28.152 49.505 28.222 50.366 ;
      RECT 28.198 49.459 28.268 50.32 ;
      RECT 28.244 49.413 28.314 50.274 ;
      RECT 28.29 49.367 28.36 50.228 ;
      RECT 28.336 49.321 28.4 50.185 ;
      RECT 28.382 49.275 28.446 50.142 ;
      RECT 28.428 49.229 28.492 50.096 ;
      RECT 28.474 49.183 28.538 50.05 ;
      RECT 28.52 49.137 28.584 50.004 ;
      RECT 28.566 49.091 28.63 49.958 ;
      RECT 28.612 49.045 28.676 49.912 ;
      RECT 28.658 48.999 28.722 49.866 ;
      RECT 28.704 48.953 28.768 49.82 ;
      RECT 28.75 48.907 28.814 49.774 ;
      RECT 28.796 48.861 28.86 49.728 ;
      RECT 28.842 48.815 28.906 49.682 ;
      RECT 28.888 48.769 28.952 49.636 ;
      RECT 28.934 48.723 28.998 49.59 ;
      RECT 28.98 48.677 29.044 49.544 ;
      RECT 29.026 48.631 29.09 49.498 ;
      RECT 29.072 48.585 29.136 49.452 ;
      RECT 29.118 48.539 29.182 49.406 ;
      RECT 29.164 48.493 29.228 49.36 ;
      RECT 29.21 48.447 29.274 49.314 ;
      RECT 29.256 48.401 29.32 49.268 ;
      RECT 29.302 48.355 29.366 49.222 ;
      RECT 29.348 48.309 29.412 49.176 ;
      RECT 29.394 48.263 29.458 49.13 ;
      RECT 29.44 48.217 29.504 49.084 ;
      RECT 29.486 48.171 29.55 49.038 ;
      RECT 29.532 48.125 29.596 48.992 ;
      RECT 29.578 48.079 29.642 48.946 ;
      RECT 29.624 48.033 29.688 48.9 ;
      RECT 29.67 47.987 29.734 48.854 ;
      RECT 29.716 47.941 29.78 48.808 ;
      RECT 29.762 47.895 29.826 48.762 ;
      RECT 29.808 47.849 29.872 48.716 ;
      RECT 29.854 47.803 29.918 48.67 ;
      RECT 29.9 47.757 29.964 48.624 ;
      RECT 29.946 47.711 30.01 48.578 ;
      RECT 29.992 47.665 30.056 48.532 ;
      RECT 30.038 47.619 30.102 48.486 ;
      RECT 30.084 47.573 30.148 48.44 ;
      RECT 30.13 47.527 30.194 48.394 ;
      RECT 30.176 47.481 30.24 48.348 ;
      RECT 30.222 47.435 30.286 48.302 ;
      RECT 30.268 47.389 30.332 48.256 ;
      RECT 30.314 47.343 30.378 48.21 ;
      RECT 30.36 47.297 30.424 48.164 ;
      RECT 30.406 47.251 30.47 48.118 ;
      RECT 30.452 47.205 30.516 48.072 ;
      RECT 30.498 47.159 30.562 48.026 ;
      RECT 30.544 47.113 30.608 47.98 ;
      RECT 30.59 47.067 30.654 47.934 ;
      RECT 30.636 47.021 30.7 47.888 ;
      RECT 30.682 46.975 30.746 47.842 ;
      RECT 30.728 46.929 30.792 47.796 ;
      RECT 30.774 46.883 30.838 47.75 ;
      RECT 30.82 46.837 30.884 47.704 ;
      RECT 30.866 46.791 30.93 47.658 ;
      RECT 30.912 46.745 30.976 47.612 ;
      RECT 30.958 46.699 31.022 47.566 ;
      RECT 31.004 46.653 31.068 47.52 ;
      RECT 31.05 46.607 31.114 47.474 ;
      RECT 31.096 46.561 31.16 47.428 ;
      RECT 31.142 46.515 31.206 47.382 ;
      RECT 31.188 46.469 31.252 47.336 ;
      RECT 31.234 46.423 31.298 47.29 ;
      RECT 31.28 46.377 31.344 47.244 ;
      RECT 31.326 46.331 31.39 47.198 ;
      RECT 31.372 46.285 31.436 47.152 ;
      RECT 31.418 46.239 31.482 47.106 ;
      RECT 31.464 46.193 31.528 47.06 ;
      RECT 31.51 46.147 31.574 47.014 ;
      RECT 31.556 46.101 31.62 46.968 ;
      RECT 31.602 46.055 31.666 46.922 ;
      RECT 31.648 46.009 31.712 46.876 ;
      RECT 31.694 45.963 31.758 46.83 ;
      RECT 31.74 45.917 31.804 46.784 ;
      RECT 31.786 45.871 31.85 46.738 ;
      RECT 31.832 45.825 31.896 46.692 ;
      RECT 31.878 45.779 31.942 46.646 ;
      RECT 31.924 45.733 31.988 46.6 ;
      RECT 31.97 45.687 32.034 46.554 ;
      RECT 32.016 45.641 32.08 46.508 ;
      RECT 32.062 45.595 32.126 46.462 ;
      RECT 32.108 45.549 32.172 46.416 ;
      RECT 32.154 45.503 32.218 46.37 ;
      RECT 32.2 45.457 32.264 46.324 ;
      RECT 32.246 45.411 32.31 46.278 ;
      RECT 32.292 45.365 32.356 46.232 ;
      RECT 32.338 45.319 32.402 46.186 ;
      RECT 32.384 45.273 32.448 46.14 ;
      RECT 32.43 45.227 32.494 46.094 ;
      RECT 32.476 45.181 32.54 46.048 ;
      RECT 32.522 45.135 32.586 46.002 ;
      RECT 32.568 45.089 32.632 45.956 ;
      RECT 32.614 45.043 32.678 45.91 ;
      RECT 32.66 44.997 32.724 45.864 ;
      RECT 32.706 44.951 32.77 45.818 ;
      RECT 32.752 44.905 32.816 45.772 ;
      RECT 32.798 44.859 32.862 45.726 ;
      RECT 32.844 44.813 32.908 45.68 ;
      RECT 32.89 44.767 32.954 45.634 ;
      RECT 32.936 44.721 33 45.588 ;
      RECT 32.982 44.675 33.046 45.542 ;
      RECT 33.028 44.629 33.092 45.496 ;
      RECT 33.074 44.583 33.138 45.45 ;
      RECT 33.12 44.537 33.184 45.404 ;
      RECT 33.166 44.491 33.23 45.358 ;
      RECT 33.212 44.445 33.276 45.312 ;
      RECT 33.258 44.399 33.322 45.266 ;
      RECT 33.304 44.353 33.368 45.22 ;
      RECT 33.35 44.307 33.414 45.174 ;
      RECT 33.396 44.261 33.46 45.128 ;
      RECT 33.442 44.215 33.506 45.082 ;
      RECT 33.488 44.169 33.552 45.036 ;
      RECT 33.534 44.123 33.598 44.99 ;
      RECT 33.58 44.077 33.644 44.944 ;
      RECT 33.626 44.031 33.69 44.898 ;
      RECT 33.672 43.985 33.736 44.852 ;
      RECT 33.718 43.939 33.782 44.806 ;
      RECT 33.764 43.893 33.828 44.76 ;
      RECT 33.81 43.847 33.874 44.714 ;
      RECT 33.856 43.801 33.92 44.668 ;
      RECT 33.902 43.755 33.966 44.622 ;
      RECT 33.948 43.709 34.012 44.576 ;
      RECT 33.994 43.663 34.058 44.53 ;
      RECT 34.04 43.617 34.104 44.484 ;
      RECT 34.086 43.571 34.15 44.438 ;
      RECT 34.132 43.525 34.196 44.392 ;
      RECT 34.178 43.479 34.242 44.346 ;
      RECT 34.224 43.433 34.288 44.3 ;
      RECT 34.27 43.387 34.334 44.254 ;
      RECT 34.316 43.341 34.38 44.208 ;
      RECT 34.362 43.295 34.426 44.162 ;
      RECT 34.408 43.249 34.472 44.116 ;
      RECT 34.454 43.203 34.518 44.07 ;
      RECT 34.5 43.157 34.564 44.024 ;
      RECT 34.546 43.111 34.61 43.978 ;
      RECT 34.592 43.065 34.656 43.932 ;
      RECT 34.638 43.019 34.702 43.886 ;
      RECT 34.684 42.973 34.748 43.84 ;
      RECT 34.73 42.927 34.794 43.794 ;
      RECT 34.776 42.881 34.84 43.748 ;
      RECT 34.822 42.835 34.886 43.702 ;
      RECT 34.868 42.789 34.932 43.656 ;
      RECT 34.914 42.743 34.978 43.61 ;
      RECT 34.96 42.697 35.024 43.564 ;
      RECT 35.006 42.651 35.07 43.518 ;
      RECT 35.052 42.605 35.116 43.472 ;
      RECT 35.098 42.559 35.162 43.426 ;
      RECT 35.144 42.513 35.208 43.38 ;
      RECT 35.19 42.467 35.254 43.334 ;
      RECT 35.236 42.421 35.3 43.288 ;
      RECT 35.282 42.375 35.346 43.242 ;
      RECT 35.328 42.329 35.392 43.196 ;
      RECT 35.374 42.283 35.438 43.15 ;
      RECT 35.42 42.237 35.484 43.104 ;
      RECT 35.466 42.191 35.53 43.058 ;
      RECT 35.512 42.145 35.576 43.012 ;
      RECT 35.558 42.099 35.622 42.966 ;
      RECT 35.604 42.053 35.668 42.92 ;
      RECT 35.65 42.007 35.714 42.874 ;
      RECT 35.696 41.961 35.76 42.828 ;
      RECT 35.742 41.915 35.806 42.782 ;
      RECT 35.788 41.869 35.852 42.736 ;
      RECT 35.834 41.823 35.898 42.69 ;
      RECT 35.88 41.777 35.944 42.644 ;
      RECT 35.926 41.731 35.99 42.598 ;
      RECT 35.972 41.685 36.036 42.552 ;
      RECT 36.018 41.639 36.082 42.506 ;
      RECT 36.064 41.593 36.128 42.46 ;
      RECT 36.11 41.547 36.174 42.414 ;
      RECT 36.156 41.501 36.22 42.368 ;
      RECT 36.202 41.455 36.266 42.322 ;
      RECT 36.248 41.409 36.312 42.276 ;
      RECT 36.294 41.363 36.358 42.23 ;
      RECT 36.34 41.317 36.404 42.184 ;
      RECT 36.386 41.271 36.45 42.138 ;
      RECT 36.432 41.225 36.496 42.092 ;
      RECT 36.478 41.179 36.542 42.046 ;
      RECT 36.524 41.133 36.588 42 ;
      RECT 36.57 41.087 36.634 41.954 ;
      RECT 36.616 41.041 36.68 41.908 ;
      RECT 36.662 40.995 36.726 41.862 ;
      RECT 36.708 40.949 36.772 41.816 ;
      RECT 36.754 40.903 36.818 41.77 ;
      RECT 36.8 40.857 36.864 41.724 ;
      RECT 36.846 40.811 36.91 41.678 ;
      RECT 36.892 40.765 36.956 41.632 ;
      RECT 36.938 40.719 37.002 41.586 ;
      RECT 36.984 40.673 37.048 41.54 ;
      RECT 37.03 40.627 37.094 41.494 ;
      RECT 37.076 40.581 37.14 41.448 ;
      RECT 37.122 40.535 37.186 41.402 ;
      RECT 37.168 40.489 37.232 41.356 ;
      RECT 37.214 40.443 37.278 41.31 ;
      RECT 37.26 40.397 37.324 41.264 ;
      RECT 37.306 40.351 37.37 41.218 ;
      RECT 37.352 40.305 37.416 41.172 ;
      RECT 37.398 40.259 37.462 41.126 ;
      RECT 37.444 40.213 37.508 41.08 ;
      RECT 37.49 40.167 37.554 41.034 ;
      RECT 37.536 40.121 37.6 40.988 ;
      RECT 37.582 40.075 37.646 40.942 ;
      RECT 37.628 40.029 37.692 40.896 ;
      RECT 37.674 39.983 37.738 40.85 ;
      RECT 37.72 39.937 37.784 40.804 ;
      RECT 37.766 39.891 37.83 40.758 ;
      RECT 37.812 39.845 37.876 40.712 ;
      RECT 37.858 39.799 37.922 40.666 ;
      RECT 37.904 39.753 37.968 40.62 ;
      RECT 37.95 39.707 38.014 40.574 ;
      RECT 37.996 39.661 38.06 40.528 ;
      RECT 38.042 39.615 38.106 40.482 ;
      RECT 38.088 39.569 38.152 40.436 ;
      RECT 38.134 39.523 38.198 40.39 ;
      RECT 38.18 39.477 38.244 40.344 ;
      RECT 38.226 39.431 38.29 40.298 ;
      RECT 38.272 39.385 38.336 40.252 ;
      RECT 38.318 39.339 38.382 40.206 ;
      RECT 38.364 39.293 38.428 40.16 ;
      RECT 38.41 39.247 38.474 40.114 ;
      RECT 38.456 39.201 38.52 40.068 ;
      RECT 38.502 39.155 38.566 40.022 ;
      RECT 38.548 39.109 38.612 39.976 ;
      RECT 38.594 39.063 38.658 39.93 ;
      RECT 38.64 39.017 38.704 39.884 ;
      RECT 38.686 38.971 38.75 39.838 ;
      RECT 38.732 38.925 38.796 39.792 ;
      RECT 38.778 38.879 38.842 39.746 ;
      RECT 38.824 38.833 38.888 39.7 ;
      RECT 38.87 38.787 38.934 39.654 ;
      RECT 38.916 38.741 38.98 39.608 ;
      RECT 38.962 38.695 39.026 39.562 ;
      RECT 39.008 38.649 39.072 39.516 ;
      RECT 39.054 38.603 39.118 39.47 ;
      RECT 39.1 38.557 39.164 39.424 ;
      RECT 39.146 38.511 39.21 39.378 ;
      RECT 39.192 38.465 39.256 39.332 ;
      RECT 39.238 38.419 39.302 39.286 ;
      RECT 39.284 38.373 39.348 39.24 ;
      RECT 39.33 38.327 39.394 39.194 ;
      RECT 39.376 38.281 39.44 39.148 ;
      RECT 39.422 38.235 39.486 39.102 ;
      RECT 39.468 38.189 39.532 39.056 ;
      RECT 39.514 38.143 39.578 39.01 ;
      RECT 39.56 38.097 39.624 38.964 ;
      RECT 39.606 38.051 39.67 38.918 ;
      RECT 39.652 38.005 39.716 38.872 ;
      RECT 39.698 37.959 39.762 38.826 ;
      RECT 39.744 37.913 39.808 38.78 ;
      RECT 39.79 37.867 39.854 38.734 ;
      RECT 39.836 37.821 39.9 38.688 ;
      RECT 39.882 37.775 39.946 38.642 ;
      RECT 39.928 37.729 39.992 38.596 ;
      RECT 39.974 37.683 40.038 38.55 ;
      RECT 40.02 37.637 40.084 38.504 ;
      RECT 40.066 37.591 40.13 38.458 ;
      RECT 40.112 37.545 40.176 38.412 ;
      RECT 40.158 37.499 40.222 38.366 ;
      RECT 40.204 37.453 40.268 38.32 ;
      RECT 40.25 37.407 40.314 38.274 ;
      RECT 40.296 37.361 40.36 38.228 ;
      RECT 40.342 37.315 40.406 38.182 ;
      RECT 40.388 37.269 40.452 38.136 ;
      RECT 40.434 37.223 40.498 38.09 ;
      RECT 40.48 37.177 40.544 38.044 ;
      RECT 40.526 37.131 40.59 37.998 ;
      RECT 40.572 37.085 40.636 37.952 ;
      RECT 40.618 37.039 40.682 37.906 ;
      RECT 40.664 36.993 40.728 37.86 ;
      RECT 40.71 36.947 40.774 37.814 ;
      RECT 40.756 36.901 40.82 37.768 ;
      RECT 40.802 36.855 40.866 37.722 ;
      RECT 40.848 36.809 40.912 37.676 ;
      RECT 40.894 36.763 40.958 37.63 ;
      RECT 40.94 36.717 41.004 37.584 ;
      RECT 40.986 36.671 41.05 37.538 ;
      RECT 41.032 36.625 41.096 37.492 ;
      RECT 41.078 36.579 41.142 37.446 ;
      RECT 41.124 36.533 41.188 37.4 ;
      RECT 41.17 36.487 41.234 37.354 ;
      RECT 41.216 36.441 41.28 37.308 ;
      RECT 41.262 36.395 41.326 37.262 ;
      RECT 41.308 36.349 41.372 37.216 ;
      RECT 41.354 36.303 41.418 37.17 ;
      RECT 41.4 36.257 41.464 37.124 ;
      RECT 41.446 36.211 41.51 37.078 ;
      RECT 41.492 36.165 41.556 37.032 ;
      RECT 41.538 36.119 41.602 36.986 ;
      RECT 41.584 36.073 41.648 36.94 ;
      RECT 41.63 36.027 41.694 36.894 ;
      RECT 41.676 35.981 41.74 36.848 ;
      RECT 41.722 35.935 41.786 36.802 ;
      RECT 41.768 35.889 41.832 36.756 ;
      RECT 41.814 35.843 41.878 36.71 ;
      RECT 41.86 35.797 41.924 36.664 ;
      RECT 41.906 35.751 41.97 36.618 ;
      RECT 41.952 35.705 42.016 36.572 ;
      RECT 41.998 35.659 42.062 36.526 ;
      RECT 42.044 35.613 42.108 36.48 ;
      RECT 42.09 35.567 42.154 36.434 ;
      RECT 42.136 35.521 42.2 36.388 ;
      RECT 42.182 35.475 42.246 36.342 ;
      RECT 42.228 35.429 42.292 36.296 ;
      RECT 42.274 35.383 42.338 36.25 ;
      RECT 42.32 35.337 42.384 36.204 ;
      RECT 42.366 35.291 42.43 36.158 ;
      RECT 42.412 35.245 42.476 36.112 ;
      RECT 42.458 35.199 42.522 36.066 ;
      RECT 42.504 35.153 42.568 36.02 ;
      RECT 42.55 35.107 42.614 35.974 ;
      RECT 42.596 35.061 42.66 35.928 ;
      RECT 42.642 35.015 42.706 35.882 ;
      RECT 42.688 34.969 42.752 35.836 ;
      RECT 42.734 34.923 42.798 35.79 ;
      RECT 42.78 34.877 42.844 35.744 ;
      RECT 42.826 34.831 42.89 35.698 ;
      RECT 42.872 34.785 42.936 35.652 ;
      RECT 42.918 34.739 42.982 35.606 ;
      RECT 42.964 34.693 43.028 35.56 ;
      RECT 43.01 34.647 43.074 35.514 ;
      RECT 43.056 34.601 43.12 35.468 ;
      RECT 43.102 34.555 43.166 35.422 ;
      RECT 43.148 34.509 43.212 35.376 ;
      RECT 43.194 34.463 43.258 35.33 ;
      RECT 43.24 34.417 43.304 35.284 ;
      RECT 43.286 34.371 43.35 35.238 ;
      RECT 43.332 34.325 43.396 35.192 ;
      RECT 43.378 34.279 43.442 35.146 ;
      RECT 43.424 34.233 43.488 35.1 ;
      RECT 43.47 34.187 43.534 35.054 ;
      RECT 43.516 34.141 43.58 35.008 ;
      RECT 43.562 34.095 43.626 34.962 ;
      RECT 43.608 34.049 43.672 34.916 ;
      RECT 43.654 34.003 43.718 34.87 ;
      RECT 43.7 33.957 43.764 34.824 ;
      RECT 43.746 33.911 43.81 34.778 ;
      RECT 43.792 33.865 43.856 34.732 ;
      RECT 43.838 33.819 43.902 34.686 ;
      RECT 43.884 33.773 43.948 34.64 ;
      RECT 43.93 33.727 43.994 34.594 ;
      RECT 43.976 33.681 44.04 34.548 ;
      RECT 44.022 33.635 44.086 34.502 ;
      RECT 44.068 33.589 44.132 34.456 ;
      RECT 44.114 33.543 44.178 34.41 ;
      RECT 44.16 33.497 44.224 34.364 ;
      RECT 44.206 33.451 44.27 34.318 ;
      RECT 44.252 33.405 44.316 34.272 ;
      RECT 44.298 33.359 44.362 34.226 ;
      RECT 44.344 33.313 44.408 34.18 ;
      RECT 44.39 33.267 44.454 34.134 ;
      RECT 44.436 33.221 44.5 34.088 ;
      RECT 44.482 33.175 44.546 34.042 ;
      RECT 44.528 33.129 44.592 33.996 ;
      RECT 44.574 33.083 44.638 33.95 ;
      RECT 44.62 33.037 44.684 33.904 ;
      RECT 44.666 32.991 44.73 33.858 ;
      RECT 44.712 32.945 44.776 33.812 ;
      RECT 44.758 32.899 44.822 33.766 ;
      RECT 44.804 32.853 44.868 33.72 ;
      RECT 44.85 32.807 44.914 33.674 ;
      RECT 44.896 32.761 44.96 33.628 ;
      RECT 44.942 32.715 45.006 33.582 ;
      RECT 44.988 32.669 45.052 33.536 ;
      RECT 45.034 32.623 45.098 33.49 ;
      RECT 45.08 32.577 45.144 33.444 ;
      RECT 45.126 32.531 45.19 33.398 ;
      RECT 45.172 32.485 45.236 33.352 ;
      RECT 45.218 32.439 45.282 33.306 ;
      RECT 45.264 32.393 45.328 33.26 ;
      RECT 45.31 32.347 45.374 33.214 ;
      RECT 45.356 32.301 45.42 33.168 ;
      RECT 45.402 32.255 45.466 33.122 ;
      RECT 45.448 32.209 45.512 33.076 ;
      RECT 45.494 32.163 45.558 33.03 ;
      RECT 45.54 32.117 45.604 32.984 ;
      RECT 45.586 32.071 45.65 32.938 ;
      RECT 45.632 32.025 45.696 32.892 ;
      RECT 45.678 31.979 45.742 32.846 ;
      RECT 45.724 31.933 45.788 32.8 ;
      RECT 45.77 31.887 45.834 32.754 ;
      RECT 45.816 31.841 45.88 32.708 ;
      RECT 45.862 31.795 45.926 32.662 ;
      RECT 45.908 31.749 45.972 32.616 ;
      RECT 45.954 31.703 46.018 32.57 ;
      RECT 46 31.657 46.064 32.524 ;
      RECT 46.046 31.611 46.11 32.478 ;
      RECT 46.092 31.565 46.156 32.432 ;
      RECT 46.138 31.519 46.202 32.386 ;
      RECT 46.184 31.473 46.248 32.34 ;
      RECT 46.23 31.427 46.294 32.294 ;
      RECT 46.276 31.381 46.34 32.248 ;
      RECT 46.322 31.335 46.386 32.202 ;
      RECT 46.368 31.289 46.432 32.156 ;
      RECT 46.414 31.243 46.478 32.11 ;
      RECT 46.46 31.197 46.524 32.064 ;
      RECT 46.506 31.151 46.57 32.018 ;
      RECT 46.552 31.105 46.616 31.972 ;
      RECT 46.598 31.059 46.662 31.926 ;
      RECT 46.644 31.013 46.708 31.88 ;
      RECT 46.69 30.967 46.754 31.834 ;
      RECT 46.736 30.921 46.8 31.788 ;
      RECT 46.782 30.875 46.846 31.742 ;
      RECT 46.828 30.829 46.892 31.696 ;
      RECT 46.874 30.783 46.938 31.65 ;
      RECT 46.92 30.737 46.984 31.604 ;
      RECT 46.966 30.691 47.03 31.558 ;
      RECT 47.012 30.645 47.076 31.512 ;
      RECT 47.058 30.599 47.122 31.466 ;
      RECT 47.104 30.553 47.168 31.42 ;
      RECT 47.15 30.507 47.214 31.374 ;
      RECT 47.196 30.461 47.26 31.328 ;
      RECT 47.242 30.415 47.306 31.282 ;
      RECT 47.288 30.369 47.352 31.236 ;
      RECT 47.334 30.323 47.398 31.19 ;
      RECT 47.38 30.277 47.444 31.144 ;
      RECT 47.426 30.231 47.49 31.098 ;
      RECT 47.472 30.185 47.536 31.052 ;
      RECT 47.518 30.139 47.582 31.006 ;
      RECT 47.564 30.093 47.628 30.96 ;
      RECT 47.61 30.047 47.674 30.914 ;
      RECT 47.656 30.001 47.72 30.868 ;
      RECT 47.702 29.955 47.766 30.822 ;
      RECT 47.748 29.909 47.812 30.776 ;
      RECT 47.794 29.863 47.858 30.73 ;
      RECT 47.84 29.817 47.904 30.684 ;
      RECT 47.886 29.771 47.95 30.638 ;
      RECT 47.932 29.725 47.996 30.592 ;
      RECT 47.978 29.679 48.042 30.546 ;
      RECT 48.024 29.633 48.088 30.5 ;
      RECT 48.07 29.587 48.134 30.454 ;
      RECT 48.116 29.541 48.18 30.408 ;
      RECT 48.162 29.495 48.226 30.362 ;
      RECT 48.208 29.449 48.272 30.316 ;
      RECT 48.254 29.403 48.318 30.27 ;
      RECT 48.3 29.357 48.364 30.224 ;
      RECT 48.346 29.311 48.41 30.178 ;
      RECT 48.392 29.265 48.456 30.132 ;
      RECT 48.438 29.219 48.502 30.086 ;
      RECT 48.484 29.173 48.548 30.04 ;
      RECT 48.53 29.127 48.594 29.994 ;
      RECT 48.576 29.081 48.64 29.948 ;
      RECT 48.622 29.035 48.686 29.902 ;
      RECT 48.668 28.989 48.732 29.856 ;
      RECT 48.714 28.943 48.778 29.81 ;
      RECT 48.76 28.897 48.824 29.764 ;
      RECT 48.806 28.851 48.87 29.718 ;
      RECT 48.852 28.805 48.916 29.672 ;
      RECT 48.898 28.759 48.962 29.626 ;
      RECT 48.944 28.713 49.008 29.58 ;
      RECT 48.99 28.667 49.054 29.534 ;
      RECT 49.036 28.621 49.1 29.488 ;
      RECT 49.082 28.575 49.146 29.442 ;
      RECT 49.128 28.529 49.192 29.396 ;
      RECT 49.174 28.483 49.238 29.35 ;
      RECT 49.22 28.437 49.284 29.304 ;
      RECT 49.266 28.391 49.33 29.258 ;
      RECT 49.312 28.345 49.376 29.212 ;
      RECT 49.358 28.299 49.422 29.166 ;
      RECT 49.404 28.253 49.468 29.12 ;
      RECT 49.45 28.207 49.514 29.074 ;
      RECT 49.496 28.161 49.56 29.028 ;
      RECT 49.542 28.115 49.606 28.982 ;
      RECT 49.588 28.069 49.652 28.936 ;
      RECT 49.634 28.023 49.698 28.89 ;
      RECT 49.68 27.977 49.744 28.844 ;
      RECT 49.726 27.931 49.79 28.798 ;
      RECT 49.772 27.885 49.836 28.752 ;
      RECT 49.818 27.839 49.882 28.706 ;
      RECT 49.864 27.793 49.928 28.66 ;
      RECT 49.91 27.747 49.974 28.614 ;
      RECT 49.956 27.701 50.02 28.568 ;
      RECT 50.002 27.655 50.066 28.522 ;
      RECT 50.048 27.609 50.112 28.476 ;
      RECT 50.094 27.563 50.158 28.43 ;
      RECT 50.14 27.517 50.204 28.384 ;
      RECT 50.186 27.471 50.25 28.338 ;
      RECT 50.232 27.425 50.296 28.292 ;
      RECT 50.278 27.379 50.342 28.246 ;
      RECT 50.324 27.333 50.388 28.2 ;
      RECT 50.37 27.287 50.434 28.154 ;
      RECT 50.416 27.241 50.48 28.108 ;
      RECT 50.462 27.195 50.526 28.062 ;
      RECT 50.508 27.149 50.572 28.016 ;
      RECT 50.554 27.103 50.618 27.97 ;
      RECT 50.6 27.057 50.664 27.924 ;
      RECT 50.646 27.011 50.71 27.878 ;
      RECT 50.692 26.965 50.756 27.832 ;
      RECT 50.738 26.919 50.802 27.786 ;
      RECT 50.784 26.873 50.848 27.74 ;
      RECT 50.83 26.827 50.894 27.694 ;
      RECT 50.876 26.781 50.94 27.648 ;
      RECT 50.922 26.735 50.986 27.602 ;
      RECT 50.968 26.689 51.032 27.556 ;
      RECT 51.014 26.643 51.078 27.51 ;
      RECT 51.06 26.597 51.124 27.464 ;
      RECT 51.106 26.551 51.17 27.418 ;
      RECT 51.152 26.505 51.216 27.372 ;
      RECT 51.198 26.459 51.262 27.326 ;
      RECT 51.244 26.413 51.308 27.28 ;
      RECT 51.29 26.367 51.354 27.234 ;
      RECT 51.336 26.321 51.4 27.188 ;
      RECT 51.382 26.275 51.446 27.142 ;
      RECT 51.428 26.229 51.492 27.096 ;
      RECT 51.474 26.183 51.538 27.05 ;
      RECT 51.52 26.137 51.584 27.004 ;
      RECT 51.566 26.091 51.63 26.958 ;
      RECT 51.612 26.045 51.676 26.912 ;
      RECT 51.658 25.999 51.722 26.866 ;
      RECT 51.704 25.953 51.768 26.82 ;
      RECT 51.75 25.907 51.814 26.774 ;
      RECT 51.796 25.861 51.86 26.728 ;
      RECT 51.842 25.815 51.906 26.682 ;
      RECT 51.888 25.769 51.952 26.636 ;
      RECT 51.934 25.723 51.998 26.59 ;
      RECT 51.98 25.677 52.044 26.544 ;
      RECT 52.026 25.631 52.09 26.498 ;
      RECT 52.072 25.585 52.136 26.452 ;
      RECT 52.118 25.539 52.182 26.406 ;
      RECT 52.164 25.493 52.228 26.36 ;
      RECT 52.21 25.447 52.274 26.314 ;
      RECT 52.256 25.401 52.32 26.268 ;
      RECT 52.302 25.355 52.366 26.222 ;
      RECT 52.348 25.309 52.412 26.176 ;
      RECT 52.394 25.263 52.458 26.13 ;
      RECT 52.44 25.217 52.504 26.084 ;
      RECT 52.486 25.171 52.55 26.038 ;
      RECT 52.532 25.125 52.596 25.992 ;
      RECT 52.578 25.079 52.642 25.946 ;
      RECT 52.624 25.033 52.688 25.9 ;
      RECT 52.67 24.987 52.734 25.854 ;
      RECT 52.716 24.941 52.78 25.808 ;
      RECT 52.762 24.895 52.826 25.762 ;
      RECT 52.808 24.849 52.872 25.716 ;
      RECT 52.854 24.803 52.918 25.67 ;
      RECT 52.9 24.757 52.964 25.624 ;
      RECT 52.946 24.711 53.01 25.578 ;
      RECT 52.992 24.665 53.056 25.532 ;
      RECT 53.038 24.619 53.102 25.486 ;
      RECT 53.084 24.573 53.148 25.44 ;
      RECT 53.13 24.527 53.194 25.394 ;
      RECT 53.176 24.481 53.24 25.348 ;
      RECT 53.222 24.435 53.286 25.302 ;
      RECT 53.268 24.389 53.332 25.256 ;
      RECT 53.314 24.343 53.378 25.21 ;
      RECT 53.36 24.297 53.424 25.164 ;
      RECT 53.406 24.251 53.47 25.118 ;
      RECT 53.452 24.205 53.516 25.072 ;
      RECT 53.498 24.159 53.562 25.026 ;
      RECT 53.544 24.113 53.608 24.98 ;
      RECT 53.59 24.067 53.654 24.934 ;
      RECT 53.636 24.021 53.7 24.888 ;
      RECT 53.682 23.975 53.746 24.842 ;
      RECT 53.728 23.929 53.792 24.796 ;
      RECT 53.774 23.883 53.838 24.75 ;
      RECT 53.82 23.837 53.884 24.704 ;
      RECT 53.866 23.791 53.93 24.658 ;
      RECT 53.912 23.745 53.976 24.612 ;
      RECT 53.958 23.699 54.022 24.566 ;
      RECT 54.004 23.653 54.068 24.52 ;
      RECT 54.05 23.607 54.114 24.474 ;
      RECT 54.096 23.561 54.16 24.428 ;
      RECT 54.142 23.515 54.206 24.382 ;
      RECT 54.188 23.469 54.252 24.336 ;
      RECT 54.234 23.423 54.298 24.29 ;
      RECT 54.28 23.377 54.344 24.244 ;
      RECT 54.326 23.331 54.39 24.198 ;
      RECT 54.372 23.285 54.436 24.152 ;
      RECT 54.418 23.239 54.482 24.106 ;
      RECT 54.464 23.193 54.528 24.06 ;
      RECT 54.51 23.147 54.574 24.014 ;
      RECT 54.556 23.101 54.62 23.968 ;
      RECT 54.602 23.055 54.666 23.922 ;
      RECT 54.648 23.009 54.712 23.876 ;
      RECT 54.694 22.963 54.758 23.83 ;
      RECT 54.74 22.917 54.804 23.784 ;
      RECT 54.786 22.871 54.85 23.738 ;
      RECT 54.832 22.825 54.896 23.692 ;
      RECT 54.878 22.779 54.942 23.646 ;
      RECT 54.924 22.733 54.988 23.6 ;
      RECT 54.97 22.687 55.034 23.554 ;
      RECT 55.016 22.641 55.08 23.508 ;
      RECT 55.062 22.595 55.126 23.462 ;
      RECT 55.108 22.549 55.172 23.416 ;
      RECT 55.154 22.503 55.218 23.37 ;
      RECT 55.2 22.457 55.264 23.324 ;
      RECT 55.246 22.411 55.31 23.278 ;
      RECT 55.292 22.365 55.356 23.232 ;
      RECT 55.338 22.319 55.402 23.186 ;
      RECT 55.384 22.273 55.448 23.14 ;
      RECT 55.43 22.227 55.494 23.094 ;
      RECT 55.476 22.181 55.54 23.048 ;
      RECT 55.522 22.135 55.586 23.002 ;
      RECT 55.568 22.089 55.632 22.956 ;
      RECT 55.614 22.043 55.678 22.91 ;
      RECT 55.66 21.997 55.724 22.864 ;
      RECT 55.706 21.951 55.77 22.818 ;
      RECT 55.752 21.905 55.816 22.772 ;
      RECT 55.798 21.859 55.862 22.726 ;
      RECT 55.844 21.813 55.908 22.68 ;
      RECT 55.89 21.767 55.954 22.634 ;
      RECT 55.936 21.721 56 22.588 ;
      RECT 55.982 21.675 56.046 22.542 ;
      RECT 56.028 21.629 56.092 22.496 ;
      RECT 56.074 21.583 56.138 22.45 ;
      RECT 56.12 21.537 56.184 22.404 ;
      RECT 56.166 21.491 56.23 22.358 ;
      RECT 56.212 21.445 56.276 22.312 ;
      RECT 56.258 21.399 56.322 22.266 ;
      RECT 56.304 21.353 56.368 22.22 ;
      RECT 56.35 21.307 56.414 22.174 ;
      RECT 56.396 21.261 56.46 22.128 ;
      RECT 56.442 21.215 56.506 22.082 ;
      RECT 56.488 21.169 56.552 22.036 ;
      RECT 56.534 21.123 56.598 21.99 ;
      RECT 56.58 21.083 56.644 21.944 ;
      RECT 56.615 21.042 56.69 21.898 ;
      RECT 56.661 20.996 56.736 21.852 ;
      RECT 56.707 20.95 56.782 21.806 ;
      RECT 56.753 20.904 56.828 21.76 ;
      RECT 56.799 20.858 56.874 21.714 ;
      RECT 56.845 20.812 56.92 21.668 ;
      RECT 56.891 20.766 56.966 21.622 ;
      RECT 56.937 20.72 57.012 21.576 ;
      RECT 56.983 20.674 57.058 21.53 ;
      RECT 57.029 20.628 57.104 21.484 ;
      RECT 57.075 20.582 57.15 21.438 ;
      RECT 57.121 20.536 57.196 21.392 ;
      RECT 57.167 20.49 57.242 21.346 ;
      RECT 57.213 20.444 57.288 21.3 ;
      RECT 57.259 20.398 57.334 21.254 ;
      RECT 57.305 20.352 57.38 21.208 ;
      RECT 57.351 20.306 57.426 21.162 ;
      RECT 57.397 20.26 57.472 21.116 ;
      RECT 57.443 20.214 57.518 21.07 ;
      RECT 57.489 20.168 57.564 21.024 ;
      RECT 57.535 20.122 57.61 20.978 ;
      RECT 57.581 20.076 57.656 20.932 ;
      RECT 57.627 20.03 57.702 20.886 ;
      RECT 57.673 19.984 57.748 20.84 ;
      RECT 57.719 19.938 57.794 20.794 ;
      RECT 57.765 19.892 57.84 20.748 ;
      RECT 57.811 19.846 57.886 20.702 ;
      RECT 57.857 19.8 57.932 20.656 ;
      RECT 57.903 19.754 57.978 20.61 ;
      RECT 57.949 19.708 58.024 20.564 ;
      RECT 57.995 19.662 58.07 20.518 ;
      RECT 58.041 19.616 58.116 20.472 ;
      RECT 58.087 19.57 58.162 20.426 ;
      RECT 58.133 19.524 58.208 20.38 ;
      RECT 58.179 19.478 58.254 20.334 ;
      RECT 58.225 19.432 58.3 20.288 ;
      RECT 58.271 19.386 58.346 20.242 ;
      RECT 58.317 19.34 58.392 20.196 ;
      RECT 58.363 19.294 58.438 20.15 ;
      RECT 58.409 19.248 58.484 20.104 ;
      RECT 58.455 19.202 58.53 20.058 ;
      RECT 58.501 19.156 58.576 20.012 ;
      RECT 58.547 19.11 58.622 19.966 ;
      RECT 58.593 19.064 58.668 19.92 ;
      RECT 58.639 19.018 58.714 19.874 ;
      RECT 58.685 18.972 58.76 19.828 ;
      RECT 58.731 18.926 58.806 19.782 ;
      RECT 58.777 18.88 58.852 19.736 ;
      RECT 58.823 18.834 58.898 19.69 ;
      RECT 58.869 18.788 58.944 19.644 ;
      RECT 58.915 18.742 58.99 19.598 ;
      RECT 58.961 18.696 59.036 19.552 ;
      RECT 59.007 18.65 59.082 19.506 ;
      RECT 59.053 18.604 59.128 19.46 ;
      RECT 59.099 18.558 59.174 19.414 ;
      RECT 59.145 18.512 59.22 19.368 ;
      RECT 59.191 18.466 59.266 19.322 ;
      RECT 59.237 18.42 59.312 19.276 ;
      RECT 59.283 18.374 59.358 19.23 ;
      RECT 59.329 18.328 59.404 19.184 ;
      RECT 59.375 18.282 59.45 19.138 ;
      RECT 59.421 18.236 59.496 19.092 ;
      RECT 59.467 18.19 59.542 19.046 ;
      RECT 59.513 18.144 59.588 19 ;
      RECT 59.559 18.098 59.634 18.954 ;
      RECT 59.605 18.052 59.68 18.908 ;
      RECT 59.651 18.006 59.726 18.862 ;
      RECT 59.697 17.96 59.772 18.816 ;
      RECT 59.743 17.914 59.818 18.77 ;
      RECT 59.789 17.868 59.864 18.724 ;
      RECT 59.835 17.822 59.91 18.678 ;
      RECT 59.881 17.776 59.956 18.632 ;
      RECT 59.927 17.73 60.002 18.586 ;
      RECT 59.973 17.684 60.048 18.54 ;
      RECT 60.019 17.638 60.094 18.494 ;
      RECT 60.065 17.592 60.14 18.448 ;
      RECT 60.111 17.546 60.186 18.402 ;
      RECT 60.157 17.5 60.232 18.356 ;
      RECT 60.203 17.454 60.278 18.31 ;
      RECT 60.249 17.408 60.324 18.264 ;
      RECT 60.295 17.362 60.37 18.218 ;
      RECT 60.341 17.316 60.416 18.172 ;
      RECT 60.387 17.27 60.462 18.126 ;
      RECT 60.433 17.224 60.508 18.08 ;
      RECT 60.479 17.178 60.554 18.034 ;
      RECT 60.525 17.132 60.6 17.988 ;
      RECT 60.571 17.086 60.646 17.942 ;
      RECT 60.617 17.04 60.692 17.896 ;
      RECT 60.663 16.994 60.738 17.85 ;
      RECT 60.709 16.948 60.784 17.804 ;
      RECT 60.755 16.902 60.83 17.758 ;
      RECT 60.801 16.856 60.876 17.712 ;
      RECT 60.847 16.81 60.922 17.666 ;
      RECT 60.893 16.764 60.968 17.62 ;
      RECT 60.939 16.718 61.014 17.574 ;
      RECT 60.985 16.672 61.06 17.528 ;
      RECT 61.031 16.626 61.106 17.482 ;
      RECT 61.077 16.58 61.152 17.436 ;
      RECT 61.123 16.534 61.198 17.39 ;
      RECT 61.169 16.488 61.244 17.344 ;
      RECT 61.215 16.442 61.29 17.298 ;
      RECT 61.261 16.396 61.336 17.252 ;
      RECT 61.307 16.35 61.382 17.206 ;
      RECT 61.353 16.304 61.428 17.16 ;
      RECT 61.399 16.258 61.474 17.114 ;
      RECT 61.445 16.212 61.52 17.068 ;
      RECT 61.491 16.166 61.566 17.022 ;
      RECT 61.537 16.122 61.612 16.976 ;
      RECT 61.58 16.1 61.658 16.93 ;
      RECT 61.58 16.1 61.704 16.884 ;
      RECT 61.58 16.1 61.75 16.838 ;
      RECT 61.58 16.1 61.796 16.792 ;
      RECT 61.58 16.1 61.842 16.746 ;
      RECT 61.58 16.1 61.888 16.7 ;
      RECT 61.58 16.1 61.934 16.654 ;
      RECT 61.58 16.1 61.98 16.608 ;
      RECT 61.58 16.1 62.026 16.562 ;
      RECT 61.58 16.1 62.072 16.516 ;
    LAYER RDL SPACING 2 ;
      RECT -20 -20 110 110 ;
  END
END P65_1233_CORNER

MACRO P65_1233_CUT
  CLASS PAD ;
  ORIGIN 0 20 ;
  FOREIGN P65_1233_CUT 0 -20 ;
  SIZE 65 BY 130 ;
  SYMMETRY X Y R90 ;
  SITE IOSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER MET5 ;
        RECT 0 99.5 65 107.5 ;
      LAYER MET4 ;
        RECT 0 99.5 65 107.5 ;
      LAYER MET3 ;
        RECT 0 99.5 65 107.5 ;
    END
  END VDD
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET5 ;
        RECT 35.3 30.5 65 42.5 ;
        RECT 35.276 30.512 65 42.488 ;
        RECT 35.23 30.547 65 42.453 ;
        RECT 35.184 30.593 65 42.407 ;
        RECT 35.138 30.639 65 42.361 ;
        RECT 35.092 30.685 65 42.315 ;
        RECT 35.046 30.731 65 42.269 ;
        RECT 35 30.777 65 42.223 ;
        RECT 35.3 44 65 56 ;
        RECT 35.276 44.012 65 55.988 ;
        RECT 35.23 44.047 65 55.953 ;
        RECT 35.184 44.093 65 55.907 ;
        RECT 35.138 44.139 65 55.861 ;
        RECT 35.092 44.185 65 55.815 ;
        RECT 35.046 44.231 65 55.769 ;
        RECT 35 44.277 65 55.723 ;
        RECT 35.3 57.5 65 63.5 ;
        RECT 35.276 57.512 65 63.488 ;
        RECT 35.23 57.547 65 63.453 ;
        RECT 35.184 57.593 65 63.407 ;
        RECT 35.138 57.639 65 63.361 ;
        RECT 35.092 57.685 65 63.315 ;
        RECT 35.046 57.731 65 63.269 ;
        RECT 35 57.777 65 63.223 ;
        RECT 35.3 68.5 65 77 ;
        RECT 35.276 68.512 65 76.988 ;
        RECT 35.23 68.547 65 76.953 ;
        RECT 35.184 68.593 65 76.907 ;
        RECT 35.138 68.639 65 76.861 ;
        RECT 35.092 68.685 65 76.815 ;
        RECT 35.046 68.731 65 76.769 ;
        RECT 35 68.777 65 76.723 ;
      LAYER MET4 ;
        RECT 35.3 30.5 65 42.5 ;
        RECT 35.276 30.512 65 42.488 ;
        RECT 35.23 30.547 65 42.453 ;
        RECT 35.184 30.593 65 42.407 ;
        RECT 35.138 30.639 65 42.361 ;
        RECT 35.092 30.685 65 42.315 ;
        RECT 35.046 30.731 65 42.269 ;
        RECT 35 30.777 65 42.223 ;
        RECT 35.3 44 65 56 ;
        RECT 35.276 44.012 65 55.988 ;
        RECT 35.23 44.047 65 55.953 ;
        RECT 35.184 44.093 65 55.907 ;
        RECT 35.138 44.139 65 55.861 ;
        RECT 35.092 44.185 65 55.815 ;
        RECT 35.046 44.231 65 55.769 ;
        RECT 35 44.277 65 55.723 ;
        RECT 35.3 57.5 65 63.5 ;
        RECT 35.276 57.512 65 63.488 ;
        RECT 35.23 57.547 65 63.453 ;
        RECT 35.184 57.593 65 63.407 ;
        RECT 35.138 57.639 65 63.361 ;
        RECT 35.092 57.685 65 63.315 ;
        RECT 35.046 57.731 65 63.269 ;
        RECT 35 57.777 65 63.223 ;
        RECT 35.3 68.5 65 77 ;
        RECT 35.276 68.512 65 76.988 ;
        RECT 35.23 68.547 65 76.953 ;
        RECT 35.184 68.593 65 76.907 ;
        RECT 35.138 68.639 65 76.861 ;
        RECT 35.092 68.685 65 76.815 ;
        RECT 35.046 68.731 65 76.769 ;
        RECT 35 68.777 65 76.723 ;
      LAYER MET3 ;
        RECT 35.3 30.5 65 42.5 ;
        RECT 35.276 30.512 65 42.488 ;
        RECT 35.23 30.547 65 42.453 ;
        RECT 35.184 30.593 65 42.407 ;
        RECT 35.138 30.639 65 42.361 ;
        RECT 35.092 30.685 65 42.315 ;
        RECT 35.046 30.731 65 42.269 ;
        RECT 35 30.777 65 42.223 ;
        RECT 35.3 44 65 56 ;
        RECT 35.276 44.012 65 55.988 ;
        RECT 35.23 44.047 65 55.953 ;
        RECT 35.184 44.093 65 55.907 ;
        RECT 35.138 44.139 65 55.861 ;
        RECT 35.092 44.185 65 55.815 ;
        RECT 35.046 44.231 65 55.769 ;
        RECT 35 44.277 65 55.723 ;
        RECT 35.3 57.5 65 63.5 ;
        RECT 35.276 57.512 65 63.488 ;
        RECT 35.23 57.547 65 63.453 ;
        RECT 35.184 57.593 65 63.407 ;
        RECT 35.138 57.639 65 63.361 ;
        RECT 35.092 57.685 65 63.315 ;
        RECT 35.046 57.731 65 63.269 ;
        RECT 35 57.777 65 63.223 ;
        RECT 35.3 68.5 65 77 ;
        RECT 35.276 68.512 65 76.988 ;
        RECT 35.23 68.547 65 76.953 ;
        RECT 35.184 68.593 65 76.907 ;
        RECT 35.138 68.639 65 76.861 ;
        RECT 35.092 68.685 65 76.815 ;
        RECT 35.046 68.731 65 76.769 ;
        RECT 35 68.777 65 76.723 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET5 ;
        RECT 0 30.788 30 42.212 ;
        RECT 0 30.753 29.976 42.247 ;
        RECT 0 30.707 29.93 42.293 ;
        RECT 0 30.661 29.884 42.339 ;
        RECT 0 30.615 29.838 42.385 ;
        RECT 0 30.569 29.792 42.431 ;
        RECT 0 30.523 29.746 42.477 ;
        RECT 0 30.5 29.7 42.5 ;
        RECT 0 44.288 30 55.712 ;
        RECT 0 44.253 29.976 55.747 ;
        RECT 0 44.207 29.93 55.793 ;
        RECT 0 44.161 29.884 55.839 ;
        RECT 0 44.115 29.838 55.885 ;
        RECT 0 44.069 29.792 55.931 ;
        RECT 0 44.023 29.746 55.977 ;
        RECT 0 44 29.7 56 ;
        RECT 0 57.788 30 63.212 ;
        RECT 0 57.753 29.976 63.247 ;
        RECT 0 57.707 29.93 63.293 ;
        RECT 0 57.661 29.884 63.339 ;
        RECT 0 57.615 29.838 63.385 ;
        RECT 0 57.569 29.792 63.431 ;
        RECT 0 57.523 29.746 63.477 ;
        RECT 0 57.5 29.7 63.5 ;
        RECT 0 68.788 30 76.712 ;
        RECT 0 68.753 29.976 76.747 ;
        RECT 0 68.707 29.93 76.793 ;
        RECT 0 68.661 29.884 76.839 ;
        RECT 0 68.615 29.838 76.885 ;
        RECT 0 68.569 29.792 76.931 ;
        RECT 0 68.523 29.746 76.977 ;
        RECT 0 68.5 29.7 77 ;
      LAYER MET4 ;
        RECT 0 30.788 30 42.212 ;
        RECT 0 30.753 29.976 42.247 ;
        RECT 0 30.707 29.93 42.293 ;
        RECT 0 30.661 29.884 42.339 ;
        RECT 0 30.615 29.838 42.385 ;
        RECT 0 30.569 29.792 42.431 ;
        RECT 0 30.523 29.746 42.477 ;
        RECT 0 30.5 29.7 42.5 ;
        RECT 0 44.288 30 55.712 ;
        RECT 0 44.253 29.976 55.747 ;
        RECT 0 44.207 29.93 55.793 ;
        RECT 0 44.161 29.884 55.839 ;
        RECT 0 44.115 29.838 55.885 ;
        RECT 0 44.069 29.792 55.931 ;
        RECT 0 44.023 29.746 55.977 ;
        RECT 0 44 29.7 56 ;
        RECT 0 57.788 30 63.212 ;
        RECT 0 57.753 29.976 63.247 ;
        RECT 0 57.707 29.93 63.293 ;
        RECT 0 57.661 29.884 63.339 ;
        RECT 0 57.615 29.838 63.385 ;
        RECT 0 57.569 29.792 63.431 ;
        RECT 0 57.523 29.746 63.477 ;
        RECT 0 57.5 29.7 63.5 ;
        RECT 0 68.788 30 76.712 ;
        RECT 0 68.753 29.976 76.747 ;
        RECT 0 68.707 29.93 76.793 ;
        RECT 0 68.661 29.884 76.839 ;
        RECT 0 68.615 29.838 76.885 ;
        RECT 0 68.569 29.792 76.931 ;
        RECT 0 68.523 29.746 76.977 ;
        RECT 0 68.5 29.7 77 ;
      LAYER MET3 ;
        RECT 0 30.788 30 42.212 ;
        RECT 0 30.753 29.976 42.247 ;
        RECT 0 30.707 29.93 42.293 ;
        RECT 0 30.661 29.884 42.339 ;
        RECT 0 30.615 29.838 42.385 ;
        RECT 0 30.569 29.792 42.431 ;
        RECT 0 30.523 29.746 42.477 ;
        RECT 0 30.5 29.7 42.5 ;
        RECT 0 44.288 30 55.712 ;
        RECT 0 44.253 29.976 55.747 ;
        RECT 0 44.207 29.93 55.793 ;
        RECT 0 44.161 29.884 55.839 ;
        RECT 0 44.115 29.838 55.885 ;
        RECT 0 44.069 29.792 55.931 ;
        RECT 0 44.023 29.746 55.977 ;
        RECT 0 44 29.7 56 ;
        RECT 0 57.788 30 63.212 ;
        RECT 0 57.753 29.976 63.247 ;
        RECT 0 57.707 29.93 63.293 ;
        RECT 0 57.661 29.884 63.339 ;
        RECT 0 57.615 29.838 63.385 ;
        RECT 0 57.569 29.792 63.431 ;
        RECT 0 57.523 29.746 63.477 ;
        RECT 0 57.5 29.7 63.5 ;
        RECT 0 68.788 30 76.712 ;
        RECT 0 68.753 29.976 76.747 ;
        RECT 0 68.707 29.93 76.793 ;
        RECT 0 68.661 29.884 76.839 ;
        RECT 0 68.615 29.838 76.885 ;
        RECT 0 68.569 29.792 76.931 ;
        RECT 0 68.523 29.746 76.977 ;
        RECT 0 68.5 29.7 77 ;
    END
  END VDDIO
  PIN VSS
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 6.966 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 6.966 LAYER VIA4 ;
    PORT
      LAYER MET5 ;
        RECT 0 91 65 98 ;
      LAYER MET4 ;
        RECT 0 91 65 98 ;
      LAYER MET3 ;
        RECT 0 91 65 98 ;
    END
  END VSS
  PIN VSSA
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 4.1958 LAYER VIA4 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    PORT
      LAYER MET5 ;
        RECT 35.3 3.5 65 15.5 ;
        RECT 35.276 3.512 65 15.488 ;
        RECT 35.23 3.547 65 15.453 ;
        RECT 35.184 3.593 65 15.407 ;
        RECT 35.138 3.639 65 15.361 ;
        RECT 35.092 3.685 65 15.315 ;
        RECT 35.046 3.731 65 15.269 ;
        RECT 35 3.777 65 15.223 ;
        RECT 35.3 17 65 29 ;
        RECT 35.276 17.012 65 28.988 ;
        RECT 35.23 17.047 65 28.953 ;
        RECT 35.184 17.093 65 28.907 ;
        RECT 35.138 17.139 65 28.861 ;
        RECT 35.092 17.185 65 28.815 ;
        RECT 35.046 17.231 65 28.769 ;
        RECT 35 17.277 65 28.723 ;
        RECT 35.3 78.5 65 89.5 ;
        RECT 35.276 78.512 65 89.488 ;
        RECT 35.23 78.547 65 89.453 ;
        RECT 35.184 78.593 65 89.407 ;
        RECT 35.138 78.639 65 89.361 ;
        RECT 35.092 78.685 65 89.315 ;
        RECT 35.046 78.731 65 89.269 ;
        RECT 35 78.777 65 89.223 ;
      LAYER MET4 ;
        RECT 35.3 3.5 65 15.5 ;
        RECT 35.276 3.512 65 15.488 ;
        RECT 35.23 3.547 65 15.453 ;
        RECT 35.184 3.593 65 15.407 ;
        RECT 35.138 3.639 65 15.361 ;
        RECT 35.092 3.685 65 15.315 ;
        RECT 35.046 3.731 65 15.269 ;
        RECT 35 3.777 65 15.223 ;
        RECT 35.3 17 65 29 ;
        RECT 35.276 17.012 65 28.988 ;
        RECT 35.23 17.047 65 28.953 ;
        RECT 35.184 17.093 65 28.907 ;
        RECT 35.138 17.139 65 28.861 ;
        RECT 35.092 17.185 65 28.815 ;
        RECT 35.046 17.231 65 28.769 ;
        RECT 35 17.277 65 28.723 ;
        RECT 35.3 78.5 65 89.5 ;
        RECT 35.276 78.512 65 89.488 ;
        RECT 35.23 78.547 65 89.453 ;
        RECT 35.184 78.593 65 89.407 ;
        RECT 35.138 78.639 65 89.361 ;
        RECT 35.092 78.685 65 89.315 ;
        RECT 35.046 78.731 65 89.269 ;
        RECT 35 78.777 65 89.223 ;
      LAYER MET3 ;
        RECT 35.3 3.5 65 15.5 ;
        RECT 35.276 3.512 65 15.488 ;
        RECT 35.23 3.547 65 15.453 ;
        RECT 35.184 3.593 65 15.407 ;
        RECT 35.138 3.639 65 15.361 ;
        RECT 35.092 3.685 65 15.315 ;
        RECT 35.046 3.731 65 15.269 ;
        RECT 35 3.777 65 15.223 ;
        RECT 35.3 17 65 29 ;
        RECT 35.276 17.012 65 28.988 ;
        RECT 35.23 17.047 65 28.953 ;
        RECT 35.184 17.093 65 28.907 ;
        RECT 35.138 17.139 65 28.861 ;
        RECT 35.092 17.185 65 28.815 ;
        RECT 35.046 17.231 65 28.769 ;
        RECT 35 17.277 65 28.723 ;
        RECT 35.3 78.5 65 89.5 ;
        RECT 35.276 78.512 65 89.488 ;
        RECT 35.23 78.547 65 89.453 ;
        RECT 35.184 78.593 65 89.407 ;
        RECT 35.138 78.639 65 89.361 ;
        RECT 35.092 78.685 65 89.315 ;
        RECT 35.046 78.731 65 89.269 ;
        RECT 35 78.777 65 89.223 ;
    END
  END VSSA
  PIN VSSIO
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 4.3092 LAYER VIA4 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    PORT
      LAYER MET5 ;
        RECT 0 3.788 30 15.212 ;
        RECT 0 3.753 29.976 15.247 ;
        RECT 0 3.707 29.93 15.293 ;
        RECT 0 3.661 29.884 15.339 ;
        RECT 0 3.615 29.838 15.385 ;
        RECT 0 3.569 29.792 15.431 ;
        RECT 0 3.523 29.746 15.477 ;
        RECT 0 3.5 29.7 15.5 ;
        RECT 0 17.288 30 28.712 ;
        RECT 0 17.253 29.976 28.747 ;
        RECT 0 17.207 29.93 28.793 ;
        RECT 0 17.161 29.884 28.839 ;
        RECT 0 17.115 29.838 28.885 ;
        RECT 0 17.069 29.792 28.931 ;
        RECT 0 17.023 29.746 28.977 ;
        RECT 0 17 29.7 29 ;
        RECT 0 78.788 30 89.212 ;
        RECT 0 78.753 29.976 89.247 ;
        RECT 0 78.707 29.93 89.293 ;
        RECT 0 78.661 29.884 89.339 ;
        RECT 0 78.615 29.838 89.385 ;
        RECT 0 78.569 29.792 89.431 ;
        RECT 0 78.523 29.746 89.477 ;
        RECT 0 78.5 29.7 89.5 ;
      LAYER MET4 ;
        RECT 0 3.788 30 15.212 ;
        RECT 0 3.753 29.976 15.247 ;
        RECT 0 3.707 29.93 15.293 ;
        RECT 0 3.661 29.884 15.339 ;
        RECT 0 3.615 29.838 15.385 ;
        RECT 0 3.569 29.792 15.431 ;
        RECT 0 3.523 29.746 15.477 ;
        RECT 0 3.5 29.7 15.5 ;
        RECT 0 17.288 30 28.712 ;
        RECT 0 17.253 29.976 28.747 ;
        RECT 0 17.207 29.93 28.793 ;
        RECT 0 17.161 29.884 28.839 ;
        RECT 0 17.115 29.838 28.885 ;
        RECT 0 17.069 29.792 28.931 ;
        RECT 0 17.023 29.746 28.977 ;
        RECT 0 17 29.7 29 ;
        RECT 0 78.788 30 89.212 ;
        RECT 0 78.753 29.976 89.247 ;
        RECT 0 78.707 29.93 89.293 ;
        RECT 0 78.661 29.884 89.339 ;
        RECT 0 78.615 29.838 89.385 ;
        RECT 0 78.569 29.792 89.431 ;
        RECT 0 78.523 29.746 89.477 ;
        RECT 0 78.5 29.7 89.5 ;
      LAYER MET3 ;
        RECT 0 3.788 30 15.212 ;
        RECT 0 3.753 29.976 15.247 ;
        RECT 0 3.707 29.93 15.293 ;
        RECT 0 3.661 29.884 15.339 ;
        RECT 0 3.615 29.838 15.385 ;
        RECT 0 3.569 29.792 15.431 ;
        RECT 0 3.523 29.746 15.477 ;
        RECT 0 3.5 29.7 15.5 ;
        RECT 0 17.288 30 28.712 ;
        RECT 0 17.253 29.976 28.747 ;
        RECT 0 17.207 29.93 28.793 ;
        RECT 0 17.161 29.884 28.839 ;
        RECT 0 17.115 29.838 28.885 ;
        RECT 0 17.069 29.792 28.931 ;
        RECT 0 17.023 29.746 28.977 ;
        RECT 0 17 29.7 29 ;
        RECT 0 78.788 30 89.212 ;
        RECT 0 78.753 29.976 89.247 ;
        RECT 0 78.707 29.93 89.293 ;
        RECT 0 78.661 29.884 89.339 ;
        RECT 0 78.615 29.838 89.385 ;
        RECT 0 78.569 29.792 89.431 ;
        RECT 0 78.523 29.746 89.477 ;
        RECT 0 78.5 29.7 89.5 ;
    END
  END VSSIO
  OBS
    LAYER MET1 SPACING 0.09 ;
      RECT 0 -20 65 110 ;
    LAYER MET2 SPACING 0.1 ;
      RECT 0 -20 65 110 ;
    LAYER MET3 SPACING 0.1 ;
      RECT 0 89.675 65 90.825 ;
      RECT 29.875 89.663 35.125 90.825 ;
      RECT 29.875 89.652 35.101 90.825 ;
      RECT 29.921 89.628 35.101 90.825 ;
      RECT 29.921 89.606 35.055 90.825 ;
      RECT 29.967 89.582 35.055 90.825 ;
      RECT 29.967 89.56 35.009 90.825 ;
      RECT 30.013 89.536 35.009 90.825 ;
      RECT 30.013 89.514 34.963 90.825 ;
      RECT 30.059 89.49 34.963 90.825 ;
      RECT 30.059 89.468 34.917 90.825 ;
      RECT 30.105 89.444 34.917 90.825 ;
      RECT 30.105 89.422 34.871 90.825 ;
      RECT 30.151 89.398 34.871 90.825 ;
      RECT 30.151 89.387 34.825 90.825 ;
      RECT 30.175 -20 34.825 90.825 ;
      RECT 30.151 76.887 34.825 78.613 ;
      RECT 30.151 76.898 34.871 78.602 ;
      RECT 30.105 76.922 34.871 78.578 ;
      RECT 30.105 76.944 34.917 78.556 ;
      RECT 30.059 76.968 34.917 78.532 ;
      RECT 30.059 76.99 34.963 78.51 ;
      RECT 30.013 77.014 34.963 78.486 ;
      RECT 30.013 77.036 35.009 78.464 ;
      RECT 29.967 77.06 35.009 78.44 ;
      RECT 29.967 77.082 35.055 78.418 ;
      RECT 29.921 77.106 35.055 78.394 ;
      RECT 29.921 77.128 35.101 78.372 ;
      RECT 29.875 77.152 35.101 78.348 ;
      RECT 29.875 77.163 35.125 78.337 ;
      RECT 0 77.175 65 78.325 ;
      RECT 30.151 63.387 34.825 68.613 ;
      RECT 30.151 63.398 34.871 68.602 ;
      RECT 30.105 63.422 34.871 68.578 ;
      RECT 30.105 63.444 34.917 68.556 ;
      RECT 30.059 63.468 34.917 68.532 ;
      RECT 30.059 63.49 34.963 68.51 ;
      RECT 30.013 63.514 34.963 68.486 ;
      RECT 30.013 63.536 35.009 68.464 ;
      RECT 29.967 63.56 35.009 68.44 ;
      RECT 29.967 63.582 35.055 68.418 ;
      RECT 29.921 63.606 35.055 68.394 ;
      RECT 29.921 63.628 35.101 68.372 ;
      RECT 29.875 63.652 35.101 68.348 ;
      RECT 29.875 63.663 35.125 68.337 ;
      RECT 0 63.675 65 68.325 ;
      RECT 30.151 55.887 34.825 57.613 ;
      RECT 30.151 55.898 34.871 57.602 ;
      RECT 30.105 55.922 34.871 57.578 ;
      RECT 30.105 55.944 34.917 57.556 ;
      RECT 30.059 55.968 34.917 57.532 ;
      RECT 30.059 55.99 34.963 57.51 ;
      RECT 30.013 56.014 34.963 57.486 ;
      RECT 30.013 56.036 35.009 57.464 ;
      RECT 29.967 56.06 35.009 57.44 ;
      RECT 29.967 56.082 35.055 57.418 ;
      RECT 29.921 56.106 35.055 57.394 ;
      RECT 29.921 56.128 35.101 57.372 ;
      RECT 29.875 56.152 35.101 57.348 ;
      RECT 29.875 56.163 35.125 57.337 ;
      RECT 0 56.175 65 57.325 ;
      RECT 30.151 42.387 34.825 44.113 ;
      RECT 30.151 42.398 34.871 44.102 ;
      RECT 30.105 42.422 34.871 44.078 ;
      RECT 30.105 42.444 34.917 44.056 ;
      RECT 30.059 42.468 34.917 44.032 ;
      RECT 30.059 42.49 34.963 44.01 ;
      RECT 30.013 42.514 34.963 43.986 ;
      RECT 30.013 42.536 35.009 43.964 ;
      RECT 29.967 42.56 35.009 43.94 ;
      RECT 29.967 42.582 35.055 43.918 ;
      RECT 29.921 42.606 35.055 43.894 ;
      RECT 29.921 42.628 35.101 43.872 ;
      RECT 29.875 42.652 35.101 43.848 ;
      RECT 29.875 42.663 35.125 43.837 ;
      RECT 0 42.675 65 43.825 ;
      RECT 30.151 28.887 34.825 30.613 ;
      RECT 30.151 28.898 34.871 30.602 ;
      RECT 30.105 28.922 34.871 30.578 ;
      RECT 30.105 28.944 34.917 30.556 ;
      RECT 30.059 28.968 34.917 30.532 ;
      RECT 30.059 28.99 34.963 30.51 ;
      RECT 30.013 29.014 34.963 30.486 ;
      RECT 30.013 29.036 35.009 30.464 ;
      RECT 29.967 29.06 35.009 30.44 ;
      RECT 29.967 29.082 35.055 30.418 ;
      RECT 29.921 29.106 35.055 30.394 ;
      RECT 29.921 29.128 35.101 30.372 ;
      RECT 29.875 29.152 35.101 30.348 ;
      RECT 29.875 29.163 35.125 30.337 ;
      RECT 0 29.175 65 30.325 ;
      RECT 30.151 15.387 34.825 17.113 ;
      RECT 30.151 15.398 34.871 17.102 ;
      RECT 30.105 15.422 34.871 17.078 ;
      RECT 30.105 15.444 34.917 17.056 ;
      RECT 30.059 15.468 34.917 17.032 ;
      RECT 30.059 15.49 34.963 17.01 ;
      RECT 30.013 15.514 34.963 16.986 ;
      RECT 30.013 15.536 35.009 16.964 ;
      RECT 29.967 15.56 35.009 16.94 ;
      RECT 29.967 15.582 35.055 16.918 ;
      RECT 29.921 15.606 35.055 16.894 ;
      RECT 29.921 15.628 35.101 16.872 ;
      RECT 29.875 15.652 35.101 16.848 ;
      RECT 29.875 15.663 35.125 16.837 ;
      RECT 0 15.675 65 16.825 ;
      RECT 30.151 -20 34.825 3.613 ;
      RECT 30.151 -20 34.871 3.602 ;
      RECT 30.105 -20 34.871 3.578 ;
      RECT 30.105 -20 34.917 3.556 ;
      RECT 30.059 -20 34.917 3.532 ;
      RECT 30.059 -20 34.963 3.51 ;
      RECT 30.013 -20 34.963 3.486 ;
      RECT 30.013 -20 35.009 3.464 ;
      RECT 29.967 -20 35.009 3.44 ;
      RECT 29.967 -20 35.055 3.418 ;
      RECT 29.921 -20 35.055 3.394 ;
      RECT 29.921 -20 35.101 3.372 ;
      RECT 29.875 -20 35.101 3.348 ;
      RECT 29.875 -20 35.125 3.337 ;
      RECT 0 -20 65 3.325 ;
      RECT 0 98.175 65 99.325 ;
      RECT 0 107.675 65 110 ;
    LAYER MET4 SPACING 0.1 ;
      RECT 0 89.675 65 90.825 ;
      RECT 29.875 89.663 35.125 90.825 ;
      RECT 29.875 89.652 35.101 90.825 ;
      RECT 29.921 89.628 35.101 90.825 ;
      RECT 29.921 89.606 35.055 90.825 ;
      RECT 29.967 89.582 35.055 90.825 ;
      RECT 29.967 89.56 35.009 90.825 ;
      RECT 30.013 89.536 35.009 90.825 ;
      RECT 30.013 89.514 34.963 90.825 ;
      RECT 30.059 89.49 34.963 90.825 ;
      RECT 30.059 89.468 34.917 90.825 ;
      RECT 30.105 89.444 34.917 90.825 ;
      RECT 30.105 89.422 34.871 90.825 ;
      RECT 30.151 89.398 34.871 90.825 ;
      RECT 30.151 89.387 34.825 90.825 ;
      RECT 30.175 -20 34.825 90.825 ;
      RECT 30.151 76.887 34.825 78.613 ;
      RECT 30.151 76.898 34.871 78.602 ;
      RECT 30.105 76.922 34.871 78.578 ;
      RECT 30.105 76.944 34.917 78.556 ;
      RECT 30.059 76.968 34.917 78.532 ;
      RECT 30.059 76.99 34.963 78.51 ;
      RECT 30.013 77.014 34.963 78.486 ;
      RECT 30.013 77.036 35.009 78.464 ;
      RECT 29.967 77.06 35.009 78.44 ;
      RECT 29.967 77.082 35.055 78.418 ;
      RECT 29.921 77.106 35.055 78.394 ;
      RECT 29.921 77.128 35.101 78.372 ;
      RECT 29.875 77.152 35.101 78.348 ;
      RECT 29.875 77.163 35.125 78.337 ;
      RECT 0 77.175 65 78.325 ;
      RECT 30.151 63.387 34.825 68.613 ;
      RECT 30.151 63.398 34.871 68.602 ;
      RECT 30.105 63.422 34.871 68.578 ;
      RECT 30.105 63.444 34.917 68.556 ;
      RECT 30.059 63.468 34.917 68.532 ;
      RECT 30.059 63.49 34.963 68.51 ;
      RECT 30.013 63.514 34.963 68.486 ;
      RECT 30.013 63.536 35.009 68.464 ;
      RECT 29.967 63.56 35.009 68.44 ;
      RECT 29.967 63.582 35.055 68.418 ;
      RECT 29.921 63.606 35.055 68.394 ;
      RECT 29.921 63.628 35.101 68.372 ;
      RECT 29.875 63.652 35.101 68.348 ;
      RECT 29.875 63.663 35.125 68.337 ;
      RECT 0 63.675 65 68.325 ;
      RECT 30.151 55.887 34.825 57.613 ;
      RECT 30.151 55.898 34.871 57.602 ;
      RECT 30.105 55.922 34.871 57.578 ;
      RECT 30.105 55.944 34.917 57.556 ;
      RECT 30.059 55.968 34.917 57.532 ;
      RECT 30.059 55.99 34.963 57.51 ;
      RECT 30.013 56.014 34.963 57.486 ;
      RECT 30.013 56.036 35.009 57.464 ;
      RECT 29.967 56.06 35.009 57.44 ;
      RECT 29.967 56.082 35.055 57.418 ;
      RECT 29.921 56.106 35.055 57.394 ;
      RECT 29.921 56.128 35.101 57.372 ;
      RECT 29.875 56.152 35.101 57.348 ;
      RECT 29.875 56.163 35.125 57.337 ;
      RECT 0 56.175 65 57.325 ;
      RECT 30.151 42.387 34.825 44.113 ;
      RECT 30.151 42.398 34.871 44.102 ;
      RECT 30.105 42.422 34.871 44.078 ;
      RECT 30.105 42.444 34.917 44.056 ;
      RECT 30.059 42.468 34.917 44.032 ;
      RECT 30.059 42.49 34.963 44.01 ;
      RECT 30.013 42.514 34.963 43.986 ;
      RECT 30.013 42.536 35.009 43.964 ;
      RECT 29.967 42.56 35.009 43.94 ;
      RECT 29.967 42.582 35.055 43.918 ;
      RECT 29.921 42.606 35.055 43.894 ;
      RECT 29.921 42.628 35.101 43.872 ;
      RECT 29.875 42.652 35.101 43.848 ;
      RECT 29.875 42.663 35.125 43.837 ;
      RECT 0 42.675 65 43.825 ;
      RECT 30.151 28.887 34.825 30.613 ;
      RECT 30.151 28.898 34.871 30.602 ;
      RECT 30.105 28.922 34.871 30.578 ;
      RECT 30.105 28.944 34.917 30.556 ;
      RECT 30.059 28.968 34.917 30.532 ;
      RECT 30.059 28.99 34.963 30.51 ;
      RECT 30.013 29.014 34.963 30.486 ;
      RECT 30.013 29.036 35.009 30.464 ;
      RECT 29.967 29.06 35.009 30.44 ;
      RECT 29.967 29.082 35.055 30.418 ;
      RECT 29.921 29.106 35.055 30.394 ;
      RECT 29.921 29.128 35.101 30.372 ;
      RECT 29.875 29.152 35.101 30.348 ;
      RECT 29.875 29.163 35.125 30.337 ;
      RECT 0 29.175 65 30.325 ;
      RECT 30.151 15.387 34.825 17.113 ;
      RECT 30.151 15.398 34.871 17.102 ;
      RECT 30.105 15.422 34.871 17.078 ;
      RECT 30.105 15.444 34.917 17.056 ;
      RECT 30.059 15.468 34.917 17.032 ;
      RECT 30.059 15.49 34.963 17.01 ;
      RECT 30.013 15.514 34.963 16.986 ;
      RECT 30.013 15.536 35.009 16.964 ;
      RECT 29.967 15.56 35.009 16.94 ;
      RECT 29.967 15.582 35.055 16.918 ;
      RECT 29.921 15.606 35.055 16.894 ;
      RECT 29.921 15.628 35.101 16.872 ;
      RECT 29.875 15.652 35.101 16.848 ;
      RECT 29.875 15.663 35.125 16.837 ;
      RECT 0 15.675 65 16.825 ;
      RECT 30.151 -20 34.825 3.613 ;
      RECT 30.151 -20 34.871 3.602 ;
      RECT 30.105 -20 34.871 3.578 ;
      RECT 30.105 -20 34.917 3.556 ;
      RECT 30.059 -20 34.917 3.532 ;
      RECT 30.059 -20 34.963 3.51 ;
      RECT 30.013 -20 34.963 3.486 ;
      RECT 30.013 -20 35.009 3.464 ;
      RECT 29.967 -20 35.009 3.44 ;
      RECT 29.967 -20 35.055 3.418 ;
      RECT 29.921 -20 35.055 3.394 ;
      RECT 29.921 -20 35.101 3.372 ;
      RECT 29.875 -20 35.101 3.348 ;
      RECT 29.875 -20 35.125 3.337 ;
      RECT 0 -20 65 3.325 ;
      RECT 0 98.175 65 99.325 ;
      RECT 0 107.675 65 110 ;
    LAYER MET5 SPACING 0.1 ;
      RECT 0 89.83 65 90.67 ;
      RECT 30.03 89.818 34.97 90.67 ;
      RECT 30.03 89.807 34.946 90.67 ;
      RECT 30.076 89.783 34.946 90.67 ;
      RECT 30.076 89.761 34.9 90.67 ;
      RECT 30.122 89.737 34.9 90.67 ;
      RECT 30.122 89.715 34.854 90.67 ;
      RECT 30.168 89.691 34.854 90.67 ;
      RECT 30.168 89.669 34.808 90.67 ;
      RECT 30.214 89.645 34.808 90.67 ;
      RECT 30.214 89.623 34.762 90.67 ;
      RECT 30.26 89.599 34.762 90.67 ;
      RECT 30.26 89.577 34.716 90.67 ;
      RECT 30.306 89.553 34.716 90.67 ;
      RECT 30.306 89.542 34.67 90.67 ;
      RECT 30.33 -20 34.67 90.67 ;
      RECT 30.306 77.042 34.67 78.458 ;
      RECT 30.306 77.053 34.716 78.447 ;
      RECT 30.26 77.077 34.716 78.423 ;
      RECT 30.26 77.099 34.762 78.401 ;
      RECT 30.214 77.123 34.762 78.377 ;
      RECT 30.214 77.145 34.808 78.355 ;
      RECT 30.168 77.169 34.808 78.331 ;
      RECT 30.168 77.191 34.854 78.309 ;
      RECT 30.122 77.215 34.854 78.285 ;
      RECT 30.122 77.237 34.9 78.263 ;
      RECT 30.076 77.261 34.9 78.239 ;
      RECT 30.076 77.283 34.946 78.217 ;
      RECT 30.03 77.307 34.946 78.193 ;
      RECT 30.03 77.318 34.97 78.182 ;
      RECT 0 77.33 65 78.17 ;
      RECT 30.306 63.542 34.67 68.458 ;
      RECT 30.306 63.553 34.716 68.447 ;
      RECT 30.26 63.577 34.716 68.423 ;
      RECT 30.26 63.599 34.762 68.401 ;
      RECT 30.214 63.623 34.762 68.377 ;
      RECT 30.214 63.645 34.808 68.355 ;
      RECT 30.168 63.669 34.808 68.331 ;
      RECT 30.168 63.691 34.854 68.309 ;
      RECT 30.122 63.715 34.854 68.285 ;
      RECT 30.122 63.737 34.9 68.263 ;
      RECT 30.076 63.761 34.9 68.239 ;
      RECT 30.076 63.783 34.946 68.217 ;
      RECT 30.03 63.807 34.946 68.193 ;
      RECT 30.03 63.818 34.97 68.182 ;
      RECT 0 63.83 65 68.17 ;
      RECT 30.306 56.042 34.67 57.458 ;
      RECT 30.306 56.053 34.716 57.447 ;
      RECT 30.26 56.077 34.716 57.423 ;
      RECT 30.26 56.099 34.762 57.401 ;
      RECT 30.214 56.123 34.762 57.377 ;
      RECT 30.214 56.145 34.808 57.355 ;
      RECT 30.168 56.169 34.808 57.331 ;
      RECT 30.168 56.191 34.854 57.309 ;
      RECT 30.122 56.215 34.854 57.285 ;
      RECT 30.122 56.237 34.9 57.263 ;
      RECT 30.076 56.261 34.9 57.239 ;
      RECT 30.076 56.283 34.946 57.217 ;
      RECT 30.03 56.307 34.946 57.193 ;
      RECT 30.03 56.318 34.97 57.182 ;
      RECT 0 56.33 65 57.17 ;
      RECT 30.306 42.542 34.67 43.958 ;
      RECT 30.306 42.553 34.716 43.947 ;
      RECT 30.26 42.577 34.716 43.923 ;
      RECT 30.26 42.599 34.762 43.901 ;
      RECT 30.214 42.623 34.762 43.877 ;
      RECT 30.214 42.645 34.808 43.855 ;
      RECT 30.168 42.669 34.808 43.831 ;
      RECT 30.168 42.691 34.854 43.809 ;
      RECT 30.122 42.715 34.854 43.785 ;
      RECT 30.122 42.737 34.9 43.763 ;
      RECT 30.076 42.761 34.9 43.739 ;
      RECT 30.076 42.783 34.946 43.717 ;
      RECT 30.03 42.807 34.946 43.693 ;
      RECT 30.03 42.818 34.97 43.682 ;
      RECT 0 42.83 65 43.67 ;
      RECT 30.306 29.042 34.67 30.458 ;
      RECT 30.306 29.053 34.716 30.447 ;
      RECT 30.26 29.077 34.716 30.423 ;
      RECT 30.26 29.099 34.762 30.401 ;
      RECT 30.214 29.123 34.762 30.377 ;
      RECT 30.214 29.145 34.808 30.355 ;
      RECT 30.168 29.169 34.808 30.331 ;
      RECT 30.168 29.191 34.854 30.309 ;
      RECT 30.122 29.215 34.854 30.285 ;
      RECT 30.122 29.237 34.9 30.263 ;
      RECT 30.076 29.261 34.9 30.239 ;
      RECT 30.076 29.283 34.946 30.217 ;
      RECT 30.03 29.307 34.946 30.193 ;
      RECT 30.03 29.318 34.97 30.182 ;
      RECT 0 29.33 65 30.17 ;
      RECT 30.306 15.542 34.67 16.958 ;
      RECT 30.306 15.553 34.716 16.947 ;
      RECT 30.26 15.577 34.716 16.923 ;
      RECT 30.26 15.599 34.762 16.901 ;
      RECT 30.214 15.623 34.762 16.877 ;
      RECT 30.214 15.645 34.808 16.855 ;
      RECT 30.168 15.669 34.808 16.831 ;
      RECT 30.168 15.691 34.854 16.809 ;
      RECT 30.122 15.715 34.854 16.785 ;
      RECT 30.122 15.737 34.9 16.763 ;
      RECT 30.076 15.761 34.9 16.739 ;
      RECT 30.076 15.783 34.946 16.717 ;
      RECT 30.03 15.807 34.946 16.693 ;
      RECT 30.03 15.818 34.97 16.682 ;
      RECT 0 15.83 65 16.67 ;
      RECT 30.306 -20 34.67 3.458 ;
      RECT 30.306 -20 34.716 3.447 ;
      RECT 30.26 -20 34.716 3.423 ;
      RECT 30.26 -20 34.762 3.401 ;
      RECT 30.214 -20 34.762 3.377 ;
      RECT 30.214 -20 34.808 3.355 ;
      RECT 30.168 -20 34.808 3.331 ;
      RECT 30.168 -20 34.854 3.309 ;
      RECT 30.122 -20 34.854 3.285 ;
      RECT 30.122 -20 34.9 3.263 ;
      RECT 30.076 -20 34.9 3.239 ;
      RECT 30.076 -20 34.946 3.217 ;
      RECT 30.03 -20 34.946 3.193 ;
      RECT 30.03 -20 34.97 3.182 ;
      RECT 0 -20 65 3.17 ;
      RECT 0 98.33 65 99.17 ;
      RECT 0 107.83 65 110 ;
    LAYER T4M2 SPACING 0.4 ;
      RECT 30.392 89.985 34.584 90.4 ;
      RECT 30.438 89.961 34.584 90.4 ;
      RECT 30.438 89.939 34.538 90.4 ;
      RECT 30.484 89.915 34.538 90.4 ;
      RECT 30.484 89.893 34.492 90.4 ;
      RECT 30.53 89.869 34.492 90.4 ;
      RECT 30.53 89.847 34.446 90.4 ;
      RECT 30.576 89.823 34.446 90.4 ;
      RECT 30.576 89.812 34.4 90.4 ;
      RECT 30.6 -20 34.4 90.4 ;
      RECT 30.576 77.312 34.4 78.188 ;
      RECT 30.576 77.323 34.446 78.177 ;
      RECT 30.53 77.347 34.446 78.153 ;
      RECT 30.53 77.369 34.492 78.131 ;
      RECT 30.484 77.393 34.492 78.107 ;
      RECT 30.484 77.415 34.538 78.085 ;
      RECT 30.438 77.439 34.538 78.061 ;
      RECT 30.438 77.461 34.584 78.039 ;
      RECT 30.392 77.485 34.584 78.015 ;
      RECT 30.392 77.507 34.63 77.993 ;
      RECT 30.346 77.531 34.63 77.969 ;
      RECT 30.576 63.812 34.4 68.188 ;
      RECT 30.576 63.823 34.446 68.177 ;
      RECT 30.53 63.847 34.446 68.153 ;
      RECT 30.53 63.869 34.492 68.131 ;
      RECT 30.484 63.893 34.492 68.107 ;
      RECT 30.484 63.915 34.538 68.085 ;
      RECT 30.438 63.939 34.538 68.061 ;
      RECT 30.438 63.961 34.584 68.039 ;
      RECT 30.392 63.985 34.584 68.015 ;
      RECT 30.392 64.007 34.63 67.993 ;
      RECT 30.346 64.031 34.63 67.969 ;
      RECT 30.346 64.053 34.676 67.947 ;
      RECT 30.3 64.077 34.676 67.923 ;
      RECT 30.3 64.088 34.7 67.912 ;
      RECT 0 64.1 65 67.9 ;
      RECT 30.576 56.312 34.4 57.188 ;
      RECT 30.576 56.323 34.446 57.177 ;
      RECT 30.53 56.347 34.446 57.153 ;
      RECT 30.53 56.369 34.492 57.131 ;
      RECT 30.484 56.393 34.492 57.107 ;
      RECT 30.484 56.415 34.538 57.085 ;
      RECT 30.438 56.439 34.538 57.061 ;
      RECT 30.438 56.461 34.584 57.039 ;
      RECT 30.392 56.485 34.584 57.015 ;
      RECT 30.392 56.507 34.63 56.993 ;
      RECT 30.346 56.531 34.63 56.969 ;
      RECT 30.576 42.812 34.4 43.688 ;
      RECT 30.576 42.823 34.446 43.677 ;
      RECT 30.53 42.847 34.446 43.653 ;
      RECT 30.53 42.869 34.492 43.631 ;
      RECT 30.484 42.893 34.492 43.607 ;
      RECT 30.484 42.915 34.538 43.585 ;
      RECT 30.438 42.939 34.538 43.561 ;
      RECT 30.438 42.961 34.584 43.539 ;
      RECT 30.392 42.985 34.584 43.515 ;
      RECT 30.392 43.007 34.63 43.493 ;
      RECT 30.346 43.031 34.63 43.469 ;
      RECT 30.576 29.312 34.4 30.188 ;
      RECT 30.576 29.323 34.446 30.177 ;
      RECT 30.53 29.347 34.446 30.153 ;
      RECT 30.53 29.369 34.492 30.131 ;
      RECT 30.484 29.393 34.492 30.107 ;
      RECT 30.484 29.415 34.538 30.085 ;
      RECT 30.438 29.439 34.538 30.061 ;
      RECT 30.438 29.461 34.584 30.039 ;
      RECT 30.392 29.485 34.584 30.015 ;
      RECT 30.392 29.507 34.63 29.993 ;
      RECT 30.346 29.531 34.63 29.969 ;
      RECT 30.576 15.812 34.4 16.688 ;
      RECT 30.576 15.823 34.446 16.677 ;
      RECT 30.53 15.847 34.446 16.653 ;
      RECT 30.53 15.869 34.492 16.631 ;
      RECT 30.484 15.893 34.492 16.607 ;
      RECT 30.484 15.915 34.538 16.585 ;
      RECT 30.438 15.939 34.538 16.561 ;
      RECT 30.438 15.961 34.584 16.539 ;
      RECT 30.392 15.985 34.584 16.515 ;
      RECT 30.392 16.007 34.63 16.493 ;
      RECT 30.346 16.031 34.63 16.469 ;
      RECT 30.576 -20 34.4 3.188 ;
      RECT 30.576 -20 34.446 3.177 ;
      RECT 30.53 -20 34.446 3.153 ;
      RECT 30.53 -20 34.492 3.131 ;
      RECT 30.484 -20 34.492 3.107 ;
      RECT 30.484 -20 34.538 3.085 ;
      RECT 30.438 -20 34.538 3.061 ;
      RECT 30.438 -20 34.584 3.039 ;
      RECT 30.392 -20 34.584 3.015 ;
      RECT 30.392 -20 34.63 2.993 ;
      RECT 30.346 -20 34.63 2.969 ;
      RECT 30.346 -20 34.676 2.947 ;
      RECT 30.3 -20 34.676 2.923 ;
      RECT 30.3 -20 34.7 2.912 ;
      RECT 0 -20 65 2.9 ;
      RECT 0 108.1 65 110 ;
    LAYER RDL SPACING 2 ;
      RECT 0 -20 65 110 ;
  END
END P65_1233_CUT

MACRO P65_1233_FILLER0005
  CLASS PAD ;
  ORIGIN 0 20 ;
  FOREIGN P65_1233_FILLER0005 0 -20 ;
  SIZE 0.005 BY 130 ;
  SYMMETRY X Y R90 ;
  SITE IOSite ;
END P65_1233_FILLER0005

MACRO P65_1233_FILLER001
  CLASS PAD ;
  ORIGIN 0 20 ;
  FOREIGN P65_1233_FILLER001 0 -20 ;
  SIZE 0.01 BY 130 ;
  SYMMETRY X Y R90 ;
  SITE IOSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER MET5 ;
        RECT 0 99.5 0.01 107.5 ;
      LAYER MET4 ;
        RECT 0 99.5 0.01 107.5 ;
      LAYER MET3 ;
        RECT 0 99.5 0.01 107.5 ;
      LAYER MET2 ;
        RECT 0 99.5 0.01 107.5 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET5 ;
        RECT 0 30.5 0.01 42.5 ;
        RECT 0 44 0.01 56 ;
        RECT 0 57.5 0.01 63.5 ;
        RECT 0 68.5 0.01 77 ;
      LAYER MET4 ;
        RECT 0 30.5 0.01 42.5 ;
        RECT 0 44 0.01 56 ;
        RECT 0 57.5 0.01 63.5 ;
        RECT 0 68.5 0.01 77 ;
      LAYER MET3 ;
        RECT 0 30.5 0.01 42.5 ;
        RECT 0 44 0.01 56 ;
        RECT 0 57.5 0.01 63.5 ;
        RECT 0 68.5 0.01 77 ;
      LAYER MET2 ;
        RECT 0 30.5 0.01 42.5 ;
        RECT 0 44 0.01 56 ;
        RECT 0 57.5 0.01 63.5 ;
        RECT 0 68.5 0.01 77 ;
    END
  END VDDIO
  PIN VSS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET5 ;
        RECT 0 91 0.01 98 ;
      LAYER MET4 ;
        RECT 0 91 0.01 98 ;
      LAYER MET3 ;
        RECT 0 91 0.01 98 ;
      LAYER MET2 ;
        RECT 0 91 0.01 98 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET5 ;
        RECT 0 3.5 0.01 15.5 ;
        RECT 0 17 0.01 29 ;
        RECT 0 78.5 0.01 89.5 ;
      LAYER MET4 ;
        RECT 0 3.5 0.01 15.5 ;
        RECT 0 17 0.01 29 ;
        RECT 0 78.5 0.01 89.5 ;
      LAYER MET3 ;
        RECT 0 3.5 0.01 15.5 ;
        RECT 0 17 0.01 29 ;
        RECT 0 78.5 0.01 89.5 ;
      LAYER MET2 ;
        RECT 0 3.5 0.01 15.5 ;
        RECT 0 17 0.01 29 ;
        RECT 0 78.5 0.01 89.5 ;
    END
  END VSSIO
END P65_1233_FILLER001

MACRO P65_1233_FILLER01
  CLASS PAD ;
  ORIGIN 0 20 ;
  FOREIGN P65_1233_FILLER01 0 -20 ;
  SIZE 0.1 BY 130 ;
  SYMMETRY X Y R90 ;
  SITE IOSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER MET5 ;
        RECT 0 99.5 0.1 107.5 ;
      LAYER MET4 ;
        RECT 0 99.5 0.1 107.5 ;
      LAYER MET3 ;
        RECT 0 99.5 0.1 107.5 ;
      LAYER MET2 ;
        RECT 0 99.5 0.1 107.5 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET5 ;
        RECT 0 30.5 0.1 42.5 ;
        RECT 0 44 0.1 56 ;
        RECT 0 57.5 0.1 63.5 ;
        RECT 0 68.5 0.1 77 ;
      LAYER MET4 ;
        RECT 0 30.5 0.1 42.5 ;
        RECT 0 44 0.1 56 ;
        RECT 0 57.5 0.1 63.5 ;
        RECT 0 68.5 0.1 77 ;
      LAYER MET3 ;
        RECT 0 30.5 0.1 42.5 ;
        RECT 0 44 0.1 56 ;
        RECT 0 57.5 0.1 63.5 ;
        RECT 0 68.5 0.1 77 ;
      LAYER MET2 ;
        RECT 0 30.5 0.1 42.5 ;
        RECT 0 44 0.1 56 ;
        RECT 0 57.5 0.1 63.5 ;
        RECT 0 68.5 0.1 77 ;
    END
  END VDDIO
  PIN VSS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET5 ;
        RECT 0 91 0.1 98 ;
      LAYER MET4 ;
        RECT 0 91 0.1 98 ;
      LAYER MET3 ;
        RECT 0 91 0.1 98 ;
      LAYER MET2 ;
        RECT 0 91 0.1 98 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET5 ;
        RECT 0 3.5 0.1 15.5 ;
        RECT 0 17 0.1 29 ;
        RECT 0 78.5 0.1 89.5 ;
      LAYER MET4 ;
        RECT 0 3.5 0.1 15.5 ;
        RECT 0 17 0.1 29 ;
        RECT 0 78.5 0.1 89.5 ;
      LAYER MET3 ;
        RECT 0 3.5 0.1 15.5 ;
        RECT 0 17 0.1 29 ;
        RECT 0 78.5 0.1 89.5 ;
      LAYER MET2 ;
        RECT 0 3.5 0.1 15.5 ;
        RECT 0 17 0.1 29 ;
        RECT 0 78.5 0.1 89.5 ;
    END
  END VSSIO
  OBS
    LAYER MET1 SPACING 0.09 ;
      RECT 0 -20 0.1 110 ;
    LAYER MET2 SPACING 0.1 ;
      RECT 0 -20 0.1 3.325 ;
      RECT 0 15.675 0.1 16.825 ;
      RECT 0 29.175 0.1 30.325 ;
      RECT 0 42.675 0.1 43.825 ;
      RECT 0 56.175 0.1 57.325 ;
      RECT 0 63.675 0.1 68.325 ;
      RECT 0 77.175 0.1 78.325 ;
      RECT 0 89.675 0.1 90.825 ;
      RECT 0 98.175 0.1 99.325 ;
      RECT 0 107.675 0.1 110 ;
    LAYER MET3 SPACING 0.1 ;
      RECT 0 -20 0.1 3.325 ;
      RECT 0 15.675 0.1 16.825 ;
      RECT 0 29.175 0.1 30.325 ;
      RECT 0 42.675 0.1 43.825 ;
      RECT 0 56.175 0.1 57.325 ;
      RECT 0 63.675 0.1 68.325 ;
      RECT 0 77.175 0.1 78.325 ;
      RECT 0 89.675 0.1 90.825 ;
      RECT 0 98.175 0.1 99.325 ;
      RECT 0 107.675 0.1 110 ;
    LAYER MET4 SPACING 0.1 ;
      RECT 0 -20 0.1 3.325 ;
      RECT 0 15.675 0.1 16.825 ;
      RECT 0 29.175 0.1 30.325 ;
      RECT 0 42.675 0.1 43.825 ;
      RECT 0 56.175 0.1 57.325 ;
      RECT 0 63.675 0.1 68.325 ;
      RECT 0 77.175 0.1 78.325 ;
      RECT 0 89.675 0.1 90.825 ;
      RECT 0 98.175 0.1 99.325 ;
      RECT 0 107.675 0.1 110 ;
    LAYER MET5 SPACING 0.1 ;
      RECT 0 -20 0.1 3.17 ;
      RECT 0 15.83 0.1 16.67 ;
      RECT 0 29.33 0.1 30.17 ;
      RECT 0 42.83 0.1 43.67 ;
      RECT 0 56.33 0.1 57.17 ;
      RECT 0 63.83 0.1 68.17 ;
      RECT 0 77.33 0.1 78.17 ;
      RECT 0 89.83 0.1 90.67 ;
      RECT 0 98.33 0.1 99.17 ;
      RECT 0 107.83 0.1 110 ;
  END
END P65_1233_FILLER01

MACRO P65_1233_FILLER1
  CLASS PAD ;
  ORIGIN 0 20 ;
  FOREIGN P65_1233_FILLER1 0 -20 ;
  SIZE 1 BY 130 ;
  SYMMETRY X Y R90 ;
  SITE IOSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER MET5 ;
        RECT 0 99.5 1 107.5 ;
      LAYER MET4 ;
        RECT 0 99.5 1 107.5 ;
      LAYER MET3 ;
        RECT 0 99.5 1 107.5 ;
      LAYER MET2 ;
        RECT 0 99.5 1 107.5 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET5 ;
        RECT 0 30.5 1 42.5 ;
        RECT 0 44 1 56 ;
        RECT 0 57.5 1 63.5 ;
        RECT 0 68.5 1 77 ;
      LAYER MET4 ;
        RECT 0 30.5 1 42.5 ;
        RECT 0 44 1 56 ;
        RECT 0 57.5 1 63.5 ;
        RECT 0 68.5 1 77 ;
      LAYER MET3 ;
        RECT 0 30.5 1 42.5 ;
        RECT 0 44 1 56 ;
        RECT 0 57.5 1 63.5 ;
        RECT 0 68.5 1 77 ;
      LAYER MET2 ;
        RECT 0 30.5 1 42.5 ;
        RECT 0 44 1 56 ;
        RECT 0 57.5 1 63.5 ;
        RECT 0 68.5 1 77 ;
    END
  END VDDIO
  PIN VSS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET5 ;
        RECT 0 91 1 98 ;
      LAYER MET4 ;
        RECT 0 91 1 98 ;
      LAYER MET3 ;
        RECT 0 91 1 98 ;
      LAYER MET2 ;
        RECT 0 91 1 98 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET5 ;
        RECT 0 3.5 1 15.5 ;
        RECT 0 17 1 29 ;
        RECT 0 78.5 1 89.5 ;
      LAYER MET4 ;
        RECT 0 3.5 1 15.5 ;
        RECT 0 17 1 29 ;
        RECT 0 78.5 1 89.5 ;
      LAYER MET3 ;
        RECT 0 3.5 1 15.5 ;
        RECT 0 17 1 29 ;
        RECT 0 78.5 1 89.5 ;
      LAYER MET2 ;
        RECT 0 3.5 1 15.5 ;
        RECT 0 17 1 29 ;
        RECT 0 78.5 1 89.5 ;
    END
  END VSSIO
  OBS
    LAYER MET1 SPACING 0.09 ;
      RECT 0 -20 1 110 ;
    LAYER MET2 SPACING 0.1 ;
      RECT 0 -20 1 3.325 ;
      RECT 0 15.675 1 16.825 ;
      RECT 0 29.175 1 30.325 ;
      RECT 0 42.675 1 43.825 ;
      RECT 0 56.175 1 57.325 ;
      RECT 0 63.675 1 68.325 ;
      RECT 0 77.175 1 78.325 ;
      RECT 0 89.675 1 90.825 ;
      RECT 0 98.175 1 99.325 ;
      RECT 0 107.675 1 110 ;
    LAYER MET3 SPACING 0.1 ;
      RECT 0 -20 1 3.325 ;
      RECT 0 15.675 1 16.825 ;
      RECT 0 29.175 1 30.325 ;
      RECT 0 42.675 1 43.825 ;
      RECT 0 56.175 1 57.325 ;
      RECT 0 63.675 1 68.325 ;
      RECT 0 77.175 1 78.325 ;
      RECT 0 89.675 1 90.825 ;
      RECT 0 98.175 1 99.325 ;
      RECT 0 107.675 1 110 ;
    LAYER MET4 SPACING 0.1 ;
      RECT 0 -20 1 3.325 ;
      RECT 0 15.675 1 16.825 ;
      RECT 0 29.175 1 30.325 ;
      RECT 0 42.675 1 43.825 ;
      RECT 0 56.175 1 57.325 ;
      RECT 0 63.675 1 68.325 ;
      RECT 0 77.175 1 78.325 ;
      RECT 0 89.675 1 90.825 ;
      RECT 0 98.175 1 99.325 ;
      RECT 0 107.675 1 110 ;
    LAYER MET5 SPACING 0.1 ;
      RECT 0 -20 1 3.17 ;
      RECT 0 15.83 1 16.67 ;
      RECT 0 29.33 1 30.17 ;
      RECT 0 42.83 1 43.67 ;
      RECT 0 56.33 1 57.17 ;
      RECT 0 63.83 1 68.17 ;
      RECT 0 77.33 1 78.17 ;
      RECT 0 89.83 1 90.67 ;
      RECT 0 98.33 1 99.17 ;
      RECT 0 107.83 1 110 ;
    LAYER T4M2 SPACING 0.4 ;
      RECT 0 -20 1 2.9 ;
      RECT 0 64.1 1 67.9 ;
      RECT 0 108.1 1 110 ;
  END
END P65_1233_FILLER1

MACRO P65_1233_FILLER10
  CLASS PAD ;
  ORIGIN 0 20 ;
  FOREIGN P65_1233_FILLER10 0 -20 ;
  SIZE 10 BY 130 ;
  SYMMETRY X Y R90 ;
  SITE IOSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER MET5 ;
        RECT 0 99.5 10 107.5 ;
      LAYER MET4 ;
        RECT 0 99.5 10 107.5 ;
      LAYER MET3 ;
        RECT 0 99.5 10 107.5 ;
      LAYER MET2 ;
        RECT 0 99.5 10 107.5 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET5 ;
        RECT 0 30.5 10 42.5 ;
        RECT 0 44 10 56 ;
        RECT 0 57.5 10 63.5 ;
        RECT 0 68.5 10 77 ;
      LAYER MET4 ;
        RECT 0 30.5 10 42.5 ;
        RECT 0 44 10 56 ;
        RECT 0 57.5 10 63.5 ;
        RECT 0 68.5 10 77 ;
      LAYER MET3 ;
        RECT 0 30.5 10 42.5 ;
        RECT 0 44 10 56 ;
        RECT 0 57.5 10 63.5 ;
        RECT 0 68.5 10 77 ;
      LAYER MET2 ;
        RECT 0 30.5 10 42.5 ;
        RECT 0 44 10 56 ;
        RECT 0 57.5 10 63.5 ;
        RECT 0 68.5 10 77 ;
    END
  END VDDIO
  PIN VSS
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 1.7496 LAYER VIA4 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 1.7496 LAYER VIA2 ;
    PORT
      LAYER MET5 ;
        RECT 0 91 10 98 ;
      LAYER MET4 ;
        RECT 0 91 10 98 ;
      LAYER MET3 ;
        RECT 0 91 10 98 ;
      LAYER MET2 ;
        RECT 0 91 10 98 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 2.916 LAYER VIA4 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 2.916 LAYER VIA2 ;
    PORT
      LAYER MET5 ;
        RECT 0 3.5 10 15.5 ;
        RECT 0 17 10 29 ;
        RECT 0 78.5 10 89.5 ;
      LAYER MET4 ;
        RECT 0 3.5 10 15.5 ;
        RECT 0 17 10 29 ;
        RECT 0 78.5 10 89.5 ;
      LAYER MET3 ;
        RECT 0 3.5 10 15.5 ;
        RECT 0 17 10 29 ;
        RECT 0 78.5 10 89.5 ;
      LAYER MET2 ;
        RECT 0 3.5 10 15.5 ;
        RECT 0 17 10 29 ;
        RECT 0 78.5 10 89.5 ;
    END
  END VSSIO
  OBS
    LAYER MET1 SPACING 0.09 ;
      RECT 0 -20 10 110 ;
    LAYER MET2 SPACING 0.1 ;
      RECT 0 -20 10 3.325 ;
      RECT 0 15.675 10 16.825 ;
      RECT 0 29.175 10 30.325 ;
      RECT 0 42.675 10 43.825 ;
      RECT 0 56.175 10 57.325 ;
      RECT 0 63.675 10 68.325 ;
      RECT 0 77.175 10 78.325 ;
      RECT 0 89.675 10 90.825 ;
      RECT 0 98.175 10 99.325 ;
      RECT 0 107.675 10 110 ;
    LAYER MET3 SPACING 0.1 ;
      RECT 0 -20 10 3.325 ;
      RECT 0 15.675 10 16.825 ;
      RECT 0 29.175 10 30.325 ;
      RECT 0 42.675 10 43.825 ;
      RECT 0 56.175 10 57.325 ;
      RECT 0 63.675 10 68.325 ;
      RECT 0 77.175 10 78.325 ;
      RECT 0 89.675 10 90.825 ;
      RECT 0 98.175 10 99.325 ;
      RECT 0 107.675 10 110 ;
    LAYER MET4 SPACING 0.1 ;
      RECT 0 -20 10 3.325 ;
      RECT 0 15.675 10 16.825 ;
      RECT 0 29.175 10 30.325 ;
      RECT 0 42.675 10 43.825 ;
      RECT 0 56.175 10 57.325 ;
      RECT 0 63.675 10 68.325 ;
      RECT 0 77.175 10 78.325 ;
      RECT 0 89.675 10 90.825 ;
      RECT 0 98.175 10 99.325 ;
      RECT 0 107.675 10 110 ;
    LAYER MET5 SPACING 0.1 ;
      RECT 0 -20 10 3.17 ;
      RECT 0 15.83 10 16.67 ;
      RECT 0 29.33 10 30.17 ;
      RECT 0 42.83 10 43.67 ;
      RECT 0 56.33 10 57.17 ;
      RECT 0 63.83 10 68.17 ;
      RECT 0 77.33 10 78.17 ;
      RECT 0 89.83 10 90.67 ;
      RECT 0 98.33 10 99.17 ;
      RECT 0 107.83 10 110 ;
    LAYER T4M2 SPACING 0.4 ;
      RECT 0 -20 10 2.9 ;
      RECT 0 64.1 10 67.9 ;
      RECT 0 108.1 10 110 ;
    LAYER RDL SPACING 2 ;
      RECT 0 -20 10 110 ;
  END
END P65_1233_FILLER10

MACRO P65_1233_FILLER2
  CLASS PAD ;
  ORIGIN 0 20 ;
  FOREIGN P65_1233_FILLER2 0 -20 ;
  SIZE 2 BY 130 ;
  SYMMETRY X Y R90 ;
  SITE IOSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER MET5 ;
        RECT 0 99.5 2 107.5 ;
      LAYER MET4 ;
        RECT 0 99.5 2 107.5 ;
      LAYER MET3 ;
        RECT 0 99.5 2 107.5 ;
      LAYER MET2 ;
        RECT 0 99.5 2 107.5 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET5 ;
        RECT 0 30.5 2 42.5 ;
        RECT 0 44 2 56 ;
        RECT 0 57.5 2 63.5 ;
        RECT 0 68.5 2 77 ;
      LAYER MET4 ;
        RECT 0 30.5 2 42.5 ;
        RECT 0 44 2 56 ;
        RECT 0 57.5 2 63.5 ;
        RECT 0 68.5 2 77 ;
      LAYER MET3 ;
        RECT 0 30.5 2 42.5 ;
        RECT 0 44 2 56 ;
        RECT 0 57.5 2 63.5 ;
        RECT 0 68.5 2 77 ;
      LAYER MET2 ;
        RECT 0 30.5 2 42.5 ;
        RECT 0 44 2 56 ;
        RECT 0 57.5 2 63.5 ;
        RECT 0 68.5 2 77 ;
    END
  END VDDIO
  PIN VSS
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.3888 LAYER VIA4 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 0.3888 LAYER VIA2 ;
    PORT
      LAYER MET5 ;
        RECT 0 91 2 98 ;
      LAYER MET4 ;
        RECT 0 91 2 98 ;
      LAYER MET3 ;
        RECT 0 91 2 98 ;
      LAYER MET2 ;
        RECT 0 91 2 98 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.648 LAYER VIA4 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 0.648 LAYER VIA2 ;
    PORT
      LAYER MET5 ;
        RECT 0 3.5 2 15.5 ;
        RECT 0 17 2 29 ;
        RECT 0 78.5 2 89.5 ;
      LAYER MET4 ;
        RECT 0 3.5 2 15.5 ;
        RECT 0 17 2 29 ;
        RECT 0 78.5 2 89.5 ;
      LAYER MET3 ;
        RECT 0 3.5 2 15.5 ;
        RECT 0 17 2 29 ;
        RECT 0 78.5 2 89.5 ;
      LAYER MET2 ;
        RECT 0 3.5 2 15.5 ;
        RECT 0 17 2 29 ;
        RECT 0 78.5 2 89.5 ;
    END
  END VSSIO
  OBS
    LAYER MET1 SPACING 0.09 ;
      RECT 0 -20 2 110 ;
    LAYER MET2 SPACING 0.1 ;
      RECT 0 -20 2 3.325 ;
      RECT 0 15.675 2 16.825 ;
      RECT 0 29.175 2 30.325 ;
      RECT 0 42.675 2 43.825 ;
      RECT 0 56.175 2 57.325 ;
      RECT 0 63.675 2 68.325 ;
      RECT 0 77.175 2 78.325 ;
      RECT 0 89.675 2 90.825 ;
      RECT 0 98.175 2 99.325 ;
      RECT 0 107.675 2 110 ;
    LAYER MET3 SPACING 0.1 ;
      RECT 0 -20 2 3.325 ;
      RECT 0 15.675 2 16.825 ;
      RECT 0 29.175 2 30.325 ;
      RECT 0 42.675 2 43.825 ;
      RECT 0 56.175 2 57.325 ;
      RECT 0 63.675 2 68.325 ;
      RECT 0 77.175 2 78.325 ;
      RECT 0 89.675 2 90.825 ;
      RECT 0 98.175 2 99.325 ;
      RECT 0 107.675 2 110 ;
    LAYER MET4 SPACING 0.1 ;
      RECT 0 -20 2 3.325 ;
      RECT 0 15.675 2 16.825 ;
      RECT 0 29.175 2 30.325 ;
      RECT 0 42.675 2 43.825 ;
      RECT 0 56.175 2 57.325 ;
      RECT 0 63.675 2 68.325 ;
      RECT 0 77.175 2 78.325 ;
      RECT 0 89.675 2 90.825 ;
      RECT 0 98.175 2 99.325 ;
      RECT 0 107.675 2 110 ;
    LAYER MET5 SPACING 0.1 ;
      RECT 0 -20 2 3.17 ;
      RECT 0 15.83 2 16.67 ;
      RECT 0 29.33 2 30.17 ;
      RECT 0 42.83 2 43.67 ;
      RECT 0 56.33 2 57.17 ;
      RECT 0 63.83 2 68.17 ;
      RECT 0 77.33 2 78.17 ;
      RECT 0 89.83 2 90.67 ;
      RECT 0 98.33 2 99.17 ;
      RECT 0 107.83 2 110 ;
    LAYER T4M2 SPACING 0.4 ;
      RECT 0 -20 2 2.9 ;
      RECT 0 64.1 2 67.9 ;
      RECT 0 108.1 2 110 ;
  END
END P65_1233_FILLER2

MACRO P65_1233_FILLER20
  CLASS PAD ;
  ORIGIN 0 20 ;
  FOREIGN P65_1233_FILLER20 0 -20 ;
  SIZE 20 BY 130 ;
  SYMMETRY X Y R90 ;
  SITE IOSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER MET5 ;
        RECT 0 99.5 20 107.5 ;
      LAYER MET4 ;
        RECT 0 99.5 20 107.5 ;
      LAYER MET3 ;
        RECT 0 99.5 20 107.5 ;
      LAYER MET2 ;
        RECT 0 99.5 20 107.5 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET5 ;
        RECT 0 30.5 20 42.5 ;
        RECT 0 44 20 56 ;
        RECT 0 57.5 20 63.5 ;
        RECT 0 68.5 20 77 ;
      LAYER MET4 ;
        RECT 0 30.5 20 42.5 ;
        RECT 0 44 20 56 ;
        RECT 0 57.5 20 63.5 ;
        RECT 0 68.5 20 77 ;
      LAYER MET3 ;
        RECT 0 30.5 20 42.5 ;
        RECT 0 44 20 56 ;
        RECT 0 57.5 20 63.5 ;
        RECT 0 68.5 20 77 ;
      LAYER MET2 ;
        RECT 0 30.5 20 42.5 ;
        RECT 0 44 20 56 ;
        RECT 0 57.5 20 63.5 ;
        RECT 0 68.5 20 77 ;
    END
  END VDDIO
  PIN VSS
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 3.0132 LAYER VIA4 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 3.0132 LAYER VIA2 ;
    PORT
      LAYER MET5 ;
        RECT 0 91 20 98 ;
      LAYER MET4 ;
        RECT 0 91 20 98 ;
      LAYER MET3 ;
        RECT 0 91 20 98 ;
      LAYER MET2 ;
        RECT 0 91 20 98 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 5.022 LAYER VIA4 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 5.022 LAYER VIA2 ;
    PORT
      LAYER MET5 ;
        RECT 0 3.5 20 15.5 ;
        RECT 0 17 20 29 ;
        RECT 0 78.5 20 89.5 ;
      LAYER MET4 ;
        RECT 0 3.5 20 15.5 ;
        RECT 0 17 20 29 ;
        RECT 0 78.5 20 89.5 ;
      LAYER MET3 ;
        RECT 0 3.5 20 15.5 ;
        RECT 0 17 20 29 ;
        RECT 0 78.5 20 89.5 ;
      LAYER MET2 ;
        RECT 0 3.5 20 15.5 ;
        RECT 0 17 20 29 ;
        RECT 0 78.5 20 89.5 ;
    END
  END VSSIO
  OBS
    LAYER MET1 SPACING 0.09 ;
      RECT 0 -20 20 110 ;
    LAYER MET2 SPACING 0.1 ;
      RECT 0 -20 20 3.325 ;
      RECT 0 15.675 20 16.825 ;
      RECT 0 29.175 20 30.325 ;
      RECT 0 42.675 20 43.825 ;
      RECT 0 56.175 20 57.325 ;
      RECT 0 63.675 20 68.325 ;
      RECT 0 77.175 20 78.325 ;
      RECT 0 89.675 20 90.825 ;
      RECT 0 98.175 20 99.325 ;
      RECT 0 107.675 20 110 ;
    LAYER MET3 SPACING 0.1 ;
      RECT 0 -20 20 3.325 ;
      RECT 0 15.675 20 16.825 ;
      RECT 0 29.175 20 30.325 ;
      RECT 0 42.675 20 43.825 ;
      RECT 0 56.175 20 57.325 ;
      RECT 0 63.675 20 68.325 ;
      RECT 0 77.175 20 78.325 ;
      RECT 0 89.675 20 90.825 ;
      RECT 0 98.175 20 99.325 ;
      RECT 0 107.675 20 110 ;
    LAYER MET4 SPACING 0.1 ;
      RECT 0 -20 20 3.325 ;
      RECT 0 15.675 20 16.825 ;
      RECT 0 29.175 20 30.325 ;
      RECT 0 42.675 20 43.825 ;
      RECT 0 56.175 20 57.325 ;
      RECT 0 63.675 20 68.325 ;
      RECT 0 77.175 20 78.325 ;
      RECT 0 89.675 20 90.825 ;
      RECT 0 98.175 20 99.325 ;
      RECT 0 107.675 20 110 ;
    LAYER MET5 SPACING 0.1 ;
      RECT 0 -20 20 3.17 ;
      RECT 0 15.83 20 16.67 ;
      RECT 0 29.33 20 30.17 ;
      RECT 0 42.83 20 43.67 ;
      RECT 0 56.33 20 57.17 ;
      RECT 0 63.83 20 68.17 ;
      RECT 0 77.33 20 78.17 ;
      RECT 0 89.83 20 90.67 ;
      RECT 0 98.33 20 99.17 ;
      RECT 0 107.83 20 110 ;
    LAYER T4M2 SPACING 0.4 ;
      RECT 0 -20 20 2.9 ;
      RECT 0 64.1 20 67.9 ;
      RECT 0 108.1 20 110 ;
    LAYER RDL SPACING 2 ;
      RECT 0 -20 20 110 ;
  END
END P65_1233_FILLER20

MACRO P65_1233_FILLER5
  CLASS PAD ;
  ORIGIN 0 20 ;
  FOREIGN P65_1233_FILLER5 0 -20 ;
  SIZE 5 BY 130 ;
  SYMMETRY X Y R90 ;
  SITE IOSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER MET5 ;
        RECT 0 99.5 5 107.5 ;
      LAYER MET4 ;
        RECT 0 99.5 5 107.5 ;
      LAYER MET3 ;
        RECT 0 99.5 5 107.5 ;
      LAYER MET2 ;
        RECT 0 99.5 5 107.5 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET5 ;
        RECT 0 30.5 5 42.5 ;
        RECT 0 44 5 56 ;
        RECT 0 57.5 5 63.5 ;
        RECT 0 68.5 5 77 ;
      LAYER MET4 ;
        RECT 0 30.5 5 42.5 ;
        RECT 0 44 5 56 ;
        RECT 0 57.5 5 63.5 ;
        RECT 0 68.5 5 77 ;
      LAYER MET3 ;
        RECT 0 30.5 5 42.5 ;
        RECT 0 44 5 56 ;
        RECT 0 57.5 5 63.5 ;
        RECT 0 68.5 5 77 ;
      LAYER MET2 ;
        RECT 0 30.5 5 42.5 ;
        RECT 0 44 5 56 ;
        RECT 0 57.5 5 63.5 ;
        RECT 0 68.5 5 77 ;
    END
  END VDDIO
  PIN VSS
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.7776 LAYER VIA4 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 0.7776 LAYER VIA2 ;
    PORT
      LAYER MET5 ;
        RECT 0 91 5 98 ;
      LAYER MET4 ;
        RECT 0 91 5 98 ;
      LAYER MET3 ;
        RECT 0 91 5 98 ;
      LAYER MET2 ;
        RECT 0 91 5 98 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 1.296 LAYER VIA4 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 1.296 LAYER VIA2 ;
    PORT
      LAYER MET5 ;
        RECT 0 3.5 5 15.5 ;
        RECT 0 17 5 29 ;
        RECT 0 78.5 5 89.5 ;
      LAYER MET4 ;
        RECT 0 3.5 5 15.5 ;
        RECT 0 17 5 29 ;
        RECT 0 78.5 5 89.5 ;
      LAYER MET3 ;
        RECT 0 3.5 5 15.5 ;
        RECT 0 17 5 29 ;
        RECT 0 78.5 5 89.5 ;
      LAYER MET2 ;
        RECT 0 3.5 5 15.5 ;
        RECT 0 17 5 29 ;
        RECT 0 78.5 5 89.5 ;
    END
  END VSSIO
  OBS
    LAYER MET1 SPACING 0.09 ;
      RECT 0 -20 5 110 ;
    LAYER MET2 SPACING 0.1 ;
      RECT 0 -20 5 3.325 ;
      RECT 0 15.675 5 16.825 ;
      RECT 0 29.175 5 30.325 ;
      RECT 0 42.675 5 43.825 ;
      RECT 0 56.175 5 57.325 ;
      RECT 0 63.675 5 68.325 ;
      RECT 0 77.175 5 78.325 ;
      RECT 0 89.675 5 90.825 ;
      RECT 0 98.175 5 99.325 ;
      RECT 0 107.675 5 110 ;
    LAYER MET3 SPACING 0.1 ;
      RECT 0 -20 5 3.325 ;
      RECT 0 15.675 5 16.825 ;
      RECT 0 29.175 5 30.325 ;
      RECT 0 42.675 5 43.825 ;
      RECT 0 56.175 5 57.325 ;
      RECT 0 63.675 5 68.325 ;
      RECT 0 77.175 5 78.325 ;
      RECT 0 89.675 5 90.825 ;
      RECT 0 98.175 5 99.325 ;
      RECT 0 107.675 5 110 ;
    LAYER MET4 SPACING 0.1 ;
      RECT 0 -20 5 3.325 ;
      RECT 0 15.675 5 16.825 ;
      RECT 0 29.175 5 30.325 ;
      RECT 0 42.675 5 43.825 ;
      RECT 0 56.175 5 57.325 ;
      RECT 0 63.675 5 68.325 ;
      RECT 0 77.175 5 78.325 ;
      RECT 0 89.675 5 90.825 ;
      RECT 0 98.175 5 99.325 ;
      RECT 0 107.675 5 110 ;
    LAYER MET5 SPACING 0.1 ;
      RECT 0 -20 5 3.17 ;
      RECT 0 15.83 5 16.67 ;
      RECT 0 29.33 5 30.17 ;
      RECT 0 42.83 5 43.67 ;
      RECT 0 56.33 5 57.17 ;
      RECT 0 63.83 5 68.17 ;
      RECT 0 77.33 5 78.17 ;
      RECT 0 89.83 5 90.67 ;
      RECT 0 98.33 5 99.17 ;
      RECT 0 107.83 5 110 ;
    LAYER T4M2 SPACING 0.4 ;
      RECT 0 -20 5 2.9 ;
      RECT 0 64.1 5 67.9 ;
      RECT 0 108.1 5 110 ;
    LAYER RDL SPACING 2 ;
      RECT 0 -20 5 110 ;
  END
END P65_1233_FILLER5

MACRO P65_1233_FILLER50
  CLASS PAD ;
  ORIGIN 0 20 ;
  FOREIGN P65_1233_FILLER50 0 -20 ;
  SIZE 50 BY 130 ;
  SYMMETRY X Y R90 ;
  SITE IOSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER MET5 ;
        RECT 0 99.5 50 107.5 ;
      LAYER MET4 ;
        RECT 0 99.5 50 107.5 ;
      LAYER MET3 ;
        RECT 0 99.5 50 107.5 ;
      LAYER MET2 ;
        RECT 0 99.5 50 107.5 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET5 ;
        RECT 0 30.5 50 42.5 ;
        RECT 0 44 50 56 ;
        RECT 0 57.5 50 63.5 ;
        RECT 0 68.5 50 77 ;
      LAYER MET4 ;
        RECT 0 30.5 50 42.5 ;
        RECT 0 44 50 56 ;
        RECT 0 57.5 50 63.5 ;
        RECT 0 68.5 50 77 ;
      LAYER MET3 ;
        RECT 0 30.5 50 42.5 ;
        RECT 0 44 50 56 ;
        RECT 0 57.5 50 63.5 ;
        RECT 0 68.5 50 77 ;
      LAYER MET2 ;
        RECT 0 30.5 50 42.5 ;
        RECT 0 44 50 56 ;
        RECT 0 57.5 50 63.5 ;
        RECT 0 68.5 50 77 ;
    END
  END VDDIO
  PIN VSS
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 8.748 LAYER VIA4 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 8.748 LAYER VIA2 ;
    PORT
      LAYER MET5 ;
        RECT 0 91 50 98 ;
      LAYER MET4 ;
        RECT 0 91 50 98 ;
      LAYER MET3 ;
        RECT 0 91 50 98 ;
      LAYER MET2 ;
        RECT 0 91 50 98 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 14.58 LAYER VIA4 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 14.58 LAYER VIA2 ;
    PORT
      LAYER MET5 ;
        RECT 0 3.5 50 15.5 ;
        RECT 0 17 50 29 ;
        RECT 0 78.5 50 89.5 ;
      LAYER MET4 ;
        RECT 0 3.5 50 15.5 ;
        RECT 0 17 50 29 ;
        RECT 0 78.5 50 89.5 ;
      LAYER MET3 ;
        RECT 0 3.5 50 15.5 ;
        RECT 0 17 50 29 ;
        RECT 0 78.5 50 89.5 ;
      LAYER MET2 ;
        RECT 0 3.5 50 15.5 ;
        RECT 0 17 50 29 ;
        RECT 0 78.5 50 89.5 ;
    END
  END VSSIO
  OBS
    LAYER MET1 SPACING 0.09 ;
      RECT 0 -20 50 110 ;
    LAYER MET2 SPACING 0.1 ;
      RECT 0 -20 50 3.325 ;
      RECT 0 15.675 50 16.825 ;
      RECT 0 29.175 50 30.325 ;
      RECT 0 42.675 50 43.825 ;
      RECT 0 56.175 50 57.325 ;
      RECT 0 63.675 50 68.325 ;
      RECT 0 77.175 50 78.325 ;
      RECT 0 89.675 50 90.825 ;
      RECT 0 98.175 50 99.325 ;
      RECT 0 107.675 50 110 ;
    LAYER MET3 SPACING 0.1 ;
      RECT 0 -20 50 3.325 ;
      RECT 0 15.675 50 16.825 ;
      RECT 0 29.175 50 30.325 ;
      RECT 0 42.675 50 43.825 ;
      RECT 0 56.175 50 57.325 ;
      RECT 0 63.675 50 68.325 ;
      RECT 0 77.175 50 78.325 ;
      RECT 0 89.675 50 90.825 ;
      RECT 0 98.175 50 99.325 ;
      RECT 0 107.675 50 110 ;
    LAYER MET4 SPACING 0.1 ;
      RECT 0 -20 50 3.325 ;
      RECT 0 15.675 50 16.825 ;
      RECT 0 29.175 50 30.325 ;
      RECT 0 42.675 50 43.825 ;
      RECT 0 56.175 50 57.325 ;
      RECT 0 63.675 50 68.325 ;
      RECT 0 77.175 50 78.325 ;
      RECT 0 89.675 50 90.825 ;
      RECT 0 98.175 50 99.325 ;
      RECT 0 107.675 50 110 ;
    LAYER MET5 SPACING 0.1 ;
      RECT 0 -20 50 3.17 ;
      RECT 0 15.83 50 16.67 ;
      RECT 0 29.33 50 30.17 ;
      RECT 0 42.83 50 43.67 ;
      RECT 0 56.33 50 57.17 ;
      RECT 0 63.83 50 68.17 ;
      RECT 0 77.33 50 78.17 ;
      RECT 0 89.83 50 90.67 ;
      RECT 0 98.33 50 99.17 ;
      RECT 0 107.83 50 110 ;
    LAYER T4M2 SPACING 0.4 ;
      RECT 0 -20 50 2.9 ;
      RECT 0 64.1 50 67.9 ;
      RECT 0 108.1 50 110 ;
    LAYER RDL SPACING 2 ;
      RECT 0 -20 50 110 ;
  END
END P65_1233_FILLER50

MACRO P65_1233_PAR
  CLASS PAD ;
  ORIGIN 0 20 ;
  FOREIGN P65_1233_PAR 0 -20 ;
  SIZE 65 BY 130 ;
  SYMMETRY X Y R90 ;
  SITE IOSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA2 ;
    ANTENNAPARTIALCUTAREA 3.645 LAYER VIA4 ;
    PORT
      LAYER MET5 ;
        RECT 8 109 57 110 ;
      LAYER MET4 ;
        RECT 8 109 57 110 ;
      LAYER MET3 ;
        RECT 8 109 57 110 ;
      LAYER MET2 ;
        RECT 8 98.085 57 110 ;
        RECT 45.92 89.5 57 110 ;
        RECT 8 89.5 19 110 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET2 ;
        RECT 0 99.98 6.5 107.02 ;
        RECT 0 99.937 6.46 107.063 ;
        RECT 0 99.891 6.414 107.109 ;
        RECT 0 99.845 6.368 107.155 ;
        RECT 0 99.799 6.322 107.201 ;
        RECT 0 99.753 6.276 107.247 ;
        RECT 0 99.707 6.23 107.293 ;
        RECT 0 99.661 6.184 107.339 ;
        RECT 0 99.615 6.138 107.385 ;
        RECT 0 99.569 6.092 107.431 ;
        RECT 0 99.523 6.046 107.477 ;
        RECT 0 99.5 6 107.5 ;
    END
    PORT
      CLASS CORE ;
      LAYER MET5 ;
        RECT 0 99.5 65 107.5 ;
      LAYER MET4 ;
        RECT 0 99.5 65 107.5 ;
      LAYER MET3 ;
        RECT 0 99.5 65 107.5 ;
    END
  END VDD
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET5 ;
        RECT 0 68.5 65 77 ;
        RECT 0 30.788 1.5 42.212 ;
        RECT 0 30.753 1.476 42.247 ;
        RECT 0 30.707 1.43 42.293 ;
        RECT 0 30.661 1.384 42.339 ;
        RECT 0 30.615 1.338 42.385 ;
        RECT 0 30.569 1.292 42.431 ;
        RECT 0 30.523 1.246 42.477 ;
        RECT 0 30.5 1.2 42.5 ;
        RECT 0 44.288 1.5 55.712 ;
        RECT 0 44.253 1.476 55.747 ;
        RECT 0 44.207 1.43 55.793 ;
        RECT 0 44.161 1.384 55.839 ;
        RECT 0 44.115 1.338 55.885 ;
        RECT 0 44.069 1.292 55.931 ;
        RECT 0 44.023 1.246 55.977 ;
        RECT 0 44 1.2 56 ;
        RECT 0 57.788 1.5 63.212 ;
        RECT 0 57.753 1.476 63.247 ;
        RECT 0 57.707 1.43 63.293 ;
        RECT 0 57.661 1.384 63.339 ;
        RECT 0 57.615 1.338 63.385 ;
        RECT 0 57.569 1.292 63.431 ;
        RECT 0 57.523 1.246 63.477 ;
        RECT 0 57.5 1.2 63.5 ;
      LAYER MET4 ;
        RECT 0 68.5 65 77 ;
        RECT 0 30.788 1.5 42.212 ;
        RECT 0 30.753 1.476 42.247 ;
        RECT 0 30.707 1.43 42.293 ;
        RECT 0 30.661 1.384 42.339 ;
        RECT 0 30.615 1.338 42.385 ;
        RECT 0 30.569 1.292 42.431 ;
        RECT 0 30.523 1.246 42.477 ;
        RECT 0 30.5 1.2 42.5 ;
        RECT 0 44.288 1.5 55.712 ;
        RECT 0 44.253 1.476 55.747 ;
        RECT 0 44.207 1.43 55.793 ;
        RECT 0 44.161 1.384 55.839 ;
        RECT 0 44.115 1.338 55.885 ;
        RECT 0 44.069 1.292 55.931 ;
        RECT 0 44.023 1.246 55.977 ;
        RECT 0 44 1.2 56 ;
        RECT 0 57.788 1.5 63.212 ;
        RECT 0 57.753 1.476 63.247 ;
        RECT 0 57.707 1.43 63.293 ;
        RECT 0 57.661 1.384 63.339 ;
        RECT 0 57.615 1.338 63.385 ;
        RECT 0 57.569 1.292 63.431 ;
        RECT 0 57.523 1.246 63.477 ;
        RECT 0 57.5 1.2 63.5 ;
      LAYER MET3 ;
        RECT 0 68.5 65 77 ;
        RECT 0 30.788 1.5 42.212 ;
        RECT 0 30.753 1.476 42.247 ;
        RECT 0 30.707 1.43 42.293 ;
        RECT 0 30.661 1.384 42.339 ;
        RECT 0 30.615 1.338 42.385 ;
        RECT 0 30.569 1.292 42.431 ;
        RECT 0 30.523 1.246 42.477 ;
        RECT 0 30.5 1.2 42.5 ;
        RECT 0 44.288 1.5 55.712 ;
        RECT 0 44.253 1.476 55.747 ;
        RECT 0 44.207 1.43 55.793 ;
        RECT 0 44.161 1.384 55.839 ;
        RECT 0 44.115 1.338 55.885 ;
        RECT 0 44.069 1.292 55.931 ;
        RECT 0 44.023 1.246 55.977 ;
        RECT 0 44 1.2 56 ;
        RECT 0 57.788 1.5 63.212 ;
        RECT 0 57.753 1.476 63.247 ;
        RECT 0 57.707 1.43 63.293 ;
        RECT 0 57.661 1.384 63.339 ;
        RECT 0 57.615 1.338 63.385 ;
        RECT 0 57.569 1.292 63.431 ;
        RECT 0 57.523 1.246 63.477 ;
        RECT 0 57.5 1.2 63.5 ;
      LAYER MET2 ;
        RECT 0 68.5 65 77 ;
        RECT 0 57.5 65 63.5 ;
        RECT 0 44 65 56 ;
        RECT 0 30.5 65 42.5 ;
        RECT 57.015 30.5 58.205 77 ;
        RECT 51.435 30.5 52.625 77 ;
        RECT 45.855 30.5 47.045 77 ;
        RECT 40.275 30.5 41.465 77 ;
        RECT 34.695 30.5 35.885 77 ;
        RECT 29.115 30.5 30.305 77 ;
        RECT 23.535 30.5 24.725 77 ;
        RECT 17.955 30.5 19.145 77 ;
        RECT 12.375 30.5 13.565 77 ;
        RECT 6.795 30.5 7.985 77 ;
    END
  END VDDA
  PIN VSS
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 45.25 LAYER MET2 ;
    ANTENNAPARTIALCUTAREA 6.2694 LAYER VIA4 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 1.6848 LAYER VIA2 ;
    PORT
      LAYER MET5 ;
        RECT 0 91 65 98 ;
      LAYER MET4 ;
        RECT 0 91 65 98 ;
      LAYER MET3 ;
        RECT 0 91 65 98 ;
      LAYER MET2 ;
        RECT 0 91.48 6.5 97.52 ;
        RECT 0 91.437 6.46 97.563 ;
        RECT 0 91.391 6.414 97.609 ;
        RECT 0 91.345 6.368 97.655 ;
        RECT 0 91.299 6.322 97.701 ;
        RECT 0 91.253 6.276 97.747 ;
        RECT 0 91.207 6.23 97.793 ;
        RECT 0 91.161 6.184 97.839 ;
        RECT 0 91.115 6.138 97.885 ;
        RECT 0 91.069 6.092 97.931 ;
        RECT 0 91.023 6.046 97.977 ;
        RECT 0 91 6 98 ;
    END
  END VSS
  PIN VSSA
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA2 ;
    ANTENNAPARTIALCUTAREA 9.7524 LAYER VIA4 ;
    PORT
      LAYER MET5 ;
        RECT 0 78.5 65 89.5 ;
        RECT 0 3.788 1.5 15.212 ;
        RECT 0 3.753 1.476 15.247 ;
        RECT 0 3.707 1.43 15.293 ;
        RECT 0 3.661 1.384 15.339 ;
        RECT 0 3.615 1.338 15.385 ;
        RECT 0 3.569 1.292 15.431 ;
        RECT 0 3.523 1.246 15.477 ;
        RECT 0 3.5 1.2 15.5 ;
        RECT 0 17.288 1.5 28.712 ;
        RECT 0 17.253 1.476 28.747 ;
        RECT 0 17.207 1.43 28.793 ;
        RECT 0 17.161 1.384 28.839 ;
        RECT 0 17.115 1.338 28.885 ;
        RECT 0 17.069 1.292 28.931 ;
        RECT 0 17.023 1.246 28.977 ;
        RECT 0 17 1.2 29 ;
      LAYER MET4 ;
        RECT 0 78.5 65 89.5 ;
        RECT 0 3.788 1.5 15.212 ;
        RECT 0 3.753 1.476 15.247 ;
        RECT 0 3.707 1.43 15.293 ;
        RECT 0 3.661 1.384 15.339 ;
        RECT 0 3.615 1.338 15.385 ;
        RECT 0 3.569 1.292 15.431 ;
        RECT 0 3.523 1.246 15.477 ;
        RECT 0 3.5 1.2 15.5 ;
        RECT 0 17.288 1.5 28.712 ;
        RECT 0 17.253 1.476 28.747 ;
        RECT 0 17.207 1.43 28.793 ;
        RECT 0 17.161 1.384 28.839 ;
        RECT 0 17.115 1.338 28.885 ;
        RECT 0 17.069 1.292 28.931 ;
        RECT 0 17.023 1.246 28.977 ;
        RECT 0 17 1.2 29 ;
      LAYER MET3 ;
        RECT 0 78.5 65 89.5 ;
        RECT 0 3.788 1.5 15.212 ;
        RECT 0 3.753 1.476 15.247 ;
        RECT 0 3.707 1.43 15.293 ;
        RECT 0 3.661 1.384 15.339 ;
        RECT 0 3.615 1.338 15.385 ;
        RECT 0 3.569 1.292 15.431 ;
        RECT 0 3.523 1.246 15.477 ;
        RECT 0 3.5 1.2 15.5 ;
        RECT 0 17.288 1.5 28.712 ;
        RECT 0 17.253 1.476 28.747 ;
        RECT 0 17.207 1.43 28.793 ;
        RECT 0 17.161 1.384 28.839 ;
        RECT 0 17.115 1.338 28.885 ;
        RECT 0 17.069 1.292 28.931 ;
        RECT 0 17.023 1.246 28.977 ;
        RECT 0 17 1.2 29 ;
      LAYER MET2 ;
        RECT 0 17 65 29 ;
        RECT 0 3.5 65 15.5 ;
        RECT 59.805 3.5 60.995 29 ;
        RECT 54.225 3.5 55.415 29 ;
        RECT 48.645 3.5 49.835 29 ;
        RECT 43.065 3.5 44.255 29 ;
        RECT 37.485 3.5 38.675 29 ;
        RECT 31.905 3.5 33.095 29 ;
        RECT 26.325 3.5 27.515 29 ;
        RECT 20.745 3.5 21.935 29 ;
        RECT 15.165 3.5 16.355 29 ;
        RECT 9.585 3.5 10.775 29 ;
        RECT 4.005 3.5 5.195 29 ;
        RECT 0 78.98 6.5 89.02 ;
        RECT 0 78.937 6.46 89.063 ;
        RECT 0 78.891 6.414 89.109 ;
        RECT 0 78.845 6.368 89.155 ;
        RECT 0 78.799 6.322 89.201 ;
        RECT 0 78.753 6.276 89.247 ;
        RECT 0 78.707 6.23 89.293 ;
        RECT 0 78.661 6.184 89.339 ;
        RECT 0 78.615 6.138 89.385 ;
        RECT 0 78.569 6.092 89.431 ;
        RECT 0 78.523 6.046 89.477 ;
        RECT 0 78.5 6 89.5 ;
    END
  END VSSA
  PIN PAD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER T4M2 ;
        RECT 57 0.983 62 66.017 ;
        RECT 57 0.943 61.966 66.057 ;
        RECT 57 0.897 61.92 66.103 ;
        RECT 57 0.851 61.874 66.149 ;
        RECT 57 0.805 61.828 66.195 ;
        RECT 57 0.759 61.782 66.241 ;
        RECT 57 0.713 61.736 66.287 ;
        RECT 57 0.667 61.69 66.333 ;
        RECT 57 0.621 61.644 66.379 ;
        RECT 57 0.575 61.598 66.425 ;
        RECT 57 0.529 61.552 66.471 ;
        RECT 57 0.483 61.506 66.517 ;
        RECT 57 0.437 61.46 66.563 ;
        RECT 57 0.391 61.414 66.609 ;
        RECT 57 0.345 61.368 66.655 ;
        RECT 57 0.299 61.322 66.701 ;
        RECT 57 0.253 61.276 66.747 ;
        RECT 57 0.207 61.23 66.793 ;
        RECT 57 0.161 61.184 66.839 ;
        RECT 57 0.115 61.138 66.885 ;
        RECT 57 0.069 61.092 66.931 ;
        RECT 57 0.023 61.046 66.977 ;
        RECT 4 57.5 61 67 ;
        RECT 3 43.5 62 51 ;
        RECT 3 29.5 62 37 ;
        RECT 3 15.5 62 23 ;
        RECT 4 0 61 9 ;
        RECT 43 0 50.5 67 ;
        RECT 29 0 36.5 67 ;
        RECT 15 0 22.5 67 ;
        RECT 3 0.977 8.5 66.023 ;
        RECT 3.966 0.017 8.5 66.983 ;
        RECT 3.92 0.057 8.5 66.943 ;
        RECT 3.874 0.103 8.5 66.897 ;
        RECT 3.828 0.149 8.5 66.851 ;
        RECT 3.782 0.195 8.5 66.805 ;
        RECT 3.736 0.241 8.5 66.759 ;
        RECT 3.69 0.287 8.5 66.713 ;
        RECT 3.644 0.333 8.5 66.667 ;
        RECT 3.598 0.379 8.5 66.621 ;
        RECT 3.552 0.425 8.5 66.575 ;
        RECT 3.506 0.471 8.5 66.529 ;
        RECT 3.46 0.517 8.5 66.483 ;
        RECT 3.414 0.563 8.5 66.437 ;
        RECT 3.368 0.609 8.5 66.391 ;
        RECT 3.322 0.655 8.5 66.345 ;
        RECT 3.276 0.701 8.5 66.299 ;
        RECT 3.23 0.747 8.5 66.253 ;
        RECT 3.184 0.793 8.5 66.207 ;
        RECT 3.138 0.839 8.5 66.161 ;
        RECT 3.092 0.885 8.5 66.115 ;
        RECT 3.046 0.931 8.5 66.069 ;
    END
  END PAD
  OBS
    LAYER MET1 SPACING 0.09 ;
      RECT 0 -20 65 110 ;
    LAYER MET2 SPACING 0.1 ;
      RECT 57.175 77.175 65 110 ;
      RECT 0 107.675 7.825 110 ;
      RECT 6.675 77.175 7.825 110 ;
      RECT 6.175 107.652 7.825 110 ;
      RECT 6.635 107.195 7.825 110 ;
      RECT 6.221 107.606 7.825 110 ;
      RECT 6.589 107.238 7.825 110 ;
      RECT 6.267 107.56 7.825 110 ;
      RECT 6.543 107.284 7.825 110 ;
      RECT 6.313 107.514 7.825 110 ;
      RECT 6.497 107.33 7.825 110 ;
      RECT 6.359 107.468 7.825 110 ;
      RECT 6.451 107.376 7.825 110 ;
      RECT 6.405 107.422 7.825 110 ;
      RECT 6.635 97.695 7.825 99.805 ;
      RECT 6.589 97.738 7.825 99.762 ;
      RECT 6.543 97.784 7.825 99.716 ;
      RECT 6.497 97.83 7.825 99.67 ;
      RECT 6.451 97.876 7.825 99.624 ;
      RECT 6.405 97.922 7.825 99.578 ;
      RECT 6.359 97.968 7.825 99.532 ;
      RECT 6.313 98.014 7.825 99.486 ;
      RECT 6.267 98.06 7.825 99.44 ;
      RECT 6.221 98.106 7.825 99.394 ;
      RECT 6.175 98.152 7.825 99.348 ;
      RECT 0 98.175 7.825 99.325 ;
      RECT 19.175 77.175 45.745 97.91 ;
      RECT 6.635 89.195 7.825 91.305 ;
      RECT 6.589 89.238 7.825 91.262 ;
      RECT 6.543 89.284 7.825 91.216 ;
      RECT 6.497 89.33 7.825 91.17 ;
      RECT 6.451 89.376 7.825 91.124 ;
      RECT 6.405 89.422 7.825 91.078 ;
      RECT 6.359 89.468 7.825 91.032 ;
      RECT 6.313 89.514 7.825 90.986 ;
      RECT 6.267 89.56 7.825 90.94 ;
      RECT 6.221 89.606 7.825 90.894 ;
      RECT 6.175 89.652 7.825 90.848 ;
      RECT 0 89.675 7.825 90.825 ;
      RECT 6.675 77.175 65 89.325 ;
      RECT 6.635 77.175 65 78.805 ;
      RECT 6.589 77.175 65 78.762 ;
      RECT 6.543 77.175 65 78.716 ;
      RECT 6.497 77.175 65 78.67 ;
      RECT 6.451 77.175 65 78.624 ;
      RECT 6.405 77.175 65 78.578 ;
      RECT 6.359 77.175 65 78.532 ;
      RECT 6.313 77.175 65 78.486 ;
      RECT 6.267 77.175 65 78.44 ;
      RECT 6.221 77.175 65 78.394 ;
      RECT 6.175 77.175 65 78.348 ;
      RECT 0 77.175 65 78.325 ;
      RECT 0 -20 65 3.325 ;
      RECT 61.17 15.675 65 16.825 ;
      RECT 0 29.175 65 30.325 ;
      RECT 58.38 42.675 65 43.825 ;
      RECT 58.38 56.175 65 57.325 ;
      RECT 58.38 63.675 65 68.325 ;
      RECT 55.59 15.675 59.63 16.825 ;
      RECT 52.8 42.675 56.84 43.825 ;
      RECT 52.8 56.175 56.84 57.325 ;
      RECT 52.8 63.675 56.84 68.325 ;
      RECT 50.01 15.675 54.05 16.825 ;
      RECT 47.22 42.675 51.26 43.825 ;
      RECT 47.22 56.175 51.26 57.325 ;
      RECT 47.22 63.675 51.26 68.325 ;
      RECT 44.43 15.675 48.47 16.825 ;
      RECT 41.64 42.675 45.68 43.825 ;
      RECT 41.64 56.175 45.68 57.325 ;
      RECT 41.64 63.675 45.68 68.325 ;
      RECT 38.85 15.675 42.89 16.825 ;
      RECT 36.06 42.675 40.1 43.825 ;
      RECT 36.06 56.175 40.1 57.325 ;
      RECT 36.06 63.675 40.1 68.325 ;
      RECT 33.27 15.675 37.31 16.825 ;
      RECT 30.48 42.675 34.52 43.825 ;
      RECT 30.48 56.175 34.52 57.325 ;
      RECT 30.48 63.675 34.52 68.325 ;
      RECT 27.69 15.675 31.73 16.825 ;
      RECT 24.9 42.675 28.94 43.825 ;
      RECT 24.9 56.175 28.94 57.325 ;
      RECT 24.9 63.675 28.94 68.325 ;
      RECT 22.11 15.675 26.15 16.825 ;
      RECT 19.32 42.675 23.36 43.825 ;
      RECT 19.32 56.175 23.36 57.325 ;
      RECT 19.32 63.675 23.36 68.325 ;
      RECT 16.53 15.675 20.57 16.825 ;
      RECT 13.74 42.675 17.78 43.825 ;
      RECT 13.74 56.175 17.78 57.325 ;
      RECT 13.74 63.675 17.78 68.325 ;
      RECT 10.95 15.675 14.99 16.825 ;
      RECT 8.16 42.675 12.2 43.825 ;
      RECT 8.16 56.175 12.2 57.325 ;
      RECT 8.16 63.675 12.2 68.325 ;
      RECT 5.37 15.675 9.41 16.825 ;
      RECT 0 42.675 6.62 43.825 ;
      RECT 0 56.175 6.62 57.325 ;
      RECT 0 63.675 6.62 68.325 ;
      RECT 0 15.675 3.83 16.825 ;
    LAYER MET3 SPACING 0.1 ;
      RECT 58.37 63.665 65 68.325 ;
      RECT 52.79 57.5 56.85 68.325 ;
      RECT 47.21 57.5 51.27 68.325 ;
      RECT 41.63 57.5 45.69 68.325 ;
      RECT 36.05 57.5 40.11 68.325 ;
      RECT 30.47 -20 34.53 68.325 ;
      RECT 24.89 57.5 28.95 68.325 ;
      RECT 19.31 57.5 23.37 68.325 ;
      RECT 13.73 57.5 17.79 68.325 ;
      RECT 8.15 57.5 12.21 68.325 ;
      RECT 0 63.675 6.63 68.325 ;
      RECT 57 -20 62 67 ;
      RECT 1.375 63.665 65 67 ;
      RECT 3 57.5 62 67 ;
      RECT 43 -20 50.5 67 ;
      RECT 29 -20 36.5 67 ;
      RECT 15 -20 22.5 67 ;
      RECT 3 -20 8.5 67 ;
      RECT 57 56.165 65 57.335 ;
      RECT 41.63 56.165 51.27 57.335 ;
      RECT 24.89 56.165 40.11 57.335 ;
      RECT 13.73 56.165 23.37 57.335 ;
      RECT 1.375 56.165 12.21 57.335 ;
      RECT 0 56.175 12.21 57.325 ;
      RECT 3 43.5 62 51 ;
      RECT 57 42.665 65 43.835 ;
      RECT 0 42.675 12.21 43.825 ;
      RECT 52.79 42.665 56.85 51 ;
      RECT 41.63 42.665 51.27 51 ;
      RECT 24.89 42.665 40.11 51 ;
      RECT 13.73 42.665 23.37 51 ;
      RECT 1.375 42.665 12.21 43.835 ;
      RECT 3 29.165 62 37 ;
      RECT 1.375 29.165 65 30.335 ;
      RECT 0 29.175 65 30.325 ;
      RECT 3 15.5 62 23 ;
      RECT 1.375 15.665 65 16.835 ;
      RECT 0 15.675 65 16.825 ;
      RECT 3 -20 62 9 ;
      RECT 1.375 -20 65 3.335 ;
      RECT 0 -20 65 3.325 ;
      RECT 63.8 3.5 65 15.5 ;
      RECT 63.776 3.512 65 15.488 ;
      RECT 63.73 3.547 65 15.453 ;
      RECT 63.684 3.593 65 15.407 ;
      RECT 63.638 3.639 65 15.361 ;
      RECT 63.592 3.685 65 15.315 ;
      RECT 63.546 3.731 65 15.269 ;
      RECT 63.5 3.777 65 15.223 ;
      RECT 63.8 17 65 29 ;
      RECT 63.776 17.012 65 28.988 ;
      RECT 63.73 17.047 65 28.953 ;
      RECT 63.684 17.093 65 28.907 ;
      RECT 63.638 17.139 65 28.861 ;
      RECT 63.592 17.185 65 28.815 ;
      RECT 63.546 17.231 65 28.769 ;
      RECT 63.5 17.277 65 28.723 ;
      RECT 63.8 30.5 65 42.5 ;
      RECT 63.776 30.512 65 42.488 ;
      RECT 63.73 30.547 65 42.453 ;
      RECT 63.684 30.593 65 42.407 ;
      RECT 63.638 30.639 65 42.361 ;
      RECT 63.592 30.685 65 42.315 ;
      RECT 63.546 30.731 65 42.269 ;
      RECT 63.5 30.777 65 42.223 ;
      RECT 63.8 44 65 56 ;
      RECT 63.776 44.012 65 55.988 ;
      RECT 63.73 44.047 65 55.953 ;
      RECT 63.684 44.093 65 55.907 ;
      RECT 63.638 44.139 65 55.861 ;
      RECT 63.592 44.185 65 55.815 ;
      RECT 63.546 44.231 65 55.769 ;
      RECT 63.5 44.277 65 55.723 ;
      RECT 63.8 57.5 65 63.5 ;
      RECT 63.776 57.512 65 63.488 ;
      RECT 63.73 57.547 65 63.453 ;
      RECT 63.684 57.593 65 63.407 ;
      RECT 63.638 57.639 65 63.361 ;
      RECT 63.592 57.685 65 63.315 ;
      RECT 63.546 57.731 65 63.269 ;
      RECT 63.5 57.777 65 63.223 ;
      RECT 57.175 107.675 65 110 ;
      RECT 57.165 107.675 65 108.825 ;
      RECT 0 107.675 7.825 110 ;
      RECT 0 107.675 7.835 108.825 ;
      RECT 0 77.175 65 78.325 ;
      RECT 57.165 89.675 65 90.825 ;
      RECT 57.165 98.175 65 99.325 ;
      RECT 52.79 56.165 56.85 57.335 ;
      RECT 19.165 89.675 45.755 90.825 ;
      RECT 0 89.675 7.835 90.825 ;
      RECT 0 98.175 7.835 99.325 ;
    LAYER MET4 SPACING 0.1 ;
      RECT 0 63.675 65 68.325 ;
      RECT 1.675 -20 65 68.325 ;
      RECT 1.375 63.652 65 68.325 ;
      RECT 1.651 63.387 65 68.325 ;
      RECT 1.421 63.606 65 68.325 ;
      RECT 1.605 63.422 65 68.325 ;
      RECT 1.467 63.56 65 68.325 ;
      RECT 1.559 63.468 65 68.325 ;
      RECT 1.513 63.514 65 68.325 ;
      RECT 1.651 55.887 65 57.613 ;
      RECT 1.605 55.922 65 57.578 ;
      RECT 1.559 55.968 65 57.532 ;
      RECT 1.513 56.014 65 57.486 ;
      RECT 1.467 56.06 65 57.44 ;
      RECT 1.421 56.106 65 57.394 ;
      RECT 1.375 56.152 65 57.348 ;
      RECT 0 56.175 65 57.325 ;
      RECT 1.651 42.387 65 44.113 ;
      RECT 1.605 42.422 65 44.078 ;
      RECT 1.559 42.468 65 44.032 ;
      RECT 1.513 42.514 65 43.986 ;
      RECT 1.467 42.56 65 43.94 ;
      RECT 1.421 42.606 65 43.894 ;
      RECT 1.375 42.652 65 43.848 ;
      RECT 0 42.675 65 43.825 ;
      RECT 1.651 28.887 65 30.613 ;
      RECT 1.605 28.922 65 30.578 ;
      RECT 1.559 28.968 65 30.532 ;
      RECT 1.513 29.014 65 30.486 ;
      RECT 1.467 29.06 65 30.44 ;
      RECT 1.421 29.106 65 30.394 ;
      RECT 1.375 29.152 65 30.348 ;
      RECT 0 29.175 65 30.325 ;
      RECT 1.651 15.387 65 17.113 ;
      RECT 1.605 15.422 65 17.078 ;
      RECT 1.559 15.468 65 17.032 ;
      RECT 1.513 15.514 65 16.986 ;
      RECT 1.467 15.56 65 16.94 ;
      RECT 1.421 15.606 65 16.894 ;
      RECT 1.375 15.652 65 16.848 ;
      RECT 0 15.675 65 16.825 ;
      RECT 1.651 -20 65 3.613 ;
      RECT 1.605 -20 65 3.578 ;
      RECT 1.559 -20 65 3.532 ;
      RECT 1.513 -20 65 3.486 ;
      RECT 1.467 -20 65 3.44 ;
      RECT 1.421 -20 65 3.394 ;
      RECT 1.375 -20 65 3.348 ;
      RECT 0 -20 65 3.325 ;
      RECT 57.175 107.675 65 110 ;
      RECT 0 107.675 7.825 110 ;
      RECT 0 107.675 65 108.825 ;
      RECT 0 77.175 65 78.325 ;
      RECT 0 89.675 65 90.825 ;
      RECT 0 98.175 65 99.325 ;
    LAYER MET5 SPACING 0.1 ;
      RECT 0 63.83 65 68.17 ;
      RECT 1.83 -20 65 68.17 ;
      RECT 1.53 63.807 65 68.17 ;
      RECT 1.806 63.542 65 68.17 ;
      RECT 1.576 63.761 65 68.17 ;
      RECT 1.76 63.577 65 68.17 ;
      RECT 1.622 63.715 65 68.17 ;
      RECT 1.714 63.623 65 68.17 ;
      RECT 1.668 63.669 65 68.17 ;
      RECT 1.806 56.042 65 57.458 ;
      RECT 1.76 56.077 65 57.423 ;
      RECT 1.714 56.123 65 57.377 ;
      RECT 1.668 56.169 65 57.331 ;
      RECT 1.622 56.215 65 57.285 ;
      RECT 1.576 56.261 65 57.239 ;
      RECT 1.53 56.307 65 57.193 ;
      RECT 0 56.33 65 57.17 ;
      RECT 1.806 42.542 65 43.958 ;
      RECT 1.76 42.577 65 43.923 ;
      RECT 1.714 42.623 65 43.877 ;
      RECT 1.668 42.669 65 43.831 ;
      RECT 1.622 42.715 65 43.785 ;
      RECT 1.576 42.761 65 43.739 ;
      RECT 1.53 42.807 65 43.693 ;
      RECT 0 42.83 65 43.67 ;
      RECT 1.806 29.042 65 30.458 ;
      RECT 1.76 29.077 65 30.423 ;
      RECT 1.714 29.123 65 30.377 ;
      RECT 1.668 29.169 65 30.331 ;
      RECT 1.622 29.215 65 30.285 ;
      RECT 1.576 29.261 65 30.239 ;
      RECT 1.53 29.307 65 30.193 ;
      RECT 0 29.33 65 30.17 ;
      RECT 1.806 15.542 65 16.958 ;
      RECT 1.76 15.577 65 16.923 ;
      RECT 1.714 15.623 65 16.877 ;
      RECT 1.668 15.669 65 16.831 ;
      RECT 1.622 15.715 65 16.785 ;
      RECT 1.576 15.761 65 16.739 ;
      RECT 1.53 15.807 65 16.693 ;
      RECT 0 15.83 65 16.67 ;
      RECT 1.806 -20 65 3.458 ;
      RECT 1.76 -20 65 3.423 ;
      RECT 1.714 -20 65 3.377 ;
      RECT 1.668 -20 65 3.331 ;
      RECT 1.622 -20 65 3.285 ;
      RECT 1.576 -20 65 3.239 ;
      RECT 1.53 -20 65 3.193 ;
      RECT 0 -20 65 3.17 ;
      RECT 57.33 107.83 65 110 ;
      RECT 0 107.83 7.67 110 ;
      RECT 0 107.83 65 108.67 ;
      RECT 0 77.33 65 78.17 ;
      RECT 0 89.83 65 90.67 ;
      RECT 0 98.33 65 99.17 ;
    LAYER T4M2 SPACING 0.4 ;
      RECT 64.584 -20 65 -3.193 ;
      RECT 0 -20 0.428 -3.205 ;
      RECT 64.538 -20 65 -3.239 ;
      RECT 0 -20 0.474 -3.251 ;
      RECT 64.492 -20 65 -3.285 ;
      RECT 0 -20 0.52 -3.297 ;
      RECT 64.446 -20 65 -3.331 ;
      RECT 0 -20 0.566 -3.343 ;
      RECT 64.4 -20 65 -3.377 ;
      RECT 0 -20 0.6 -3.383 ;
      RECT 0 -20 65 -3.4 ;
      RECT 57.6 108.1 65 110 ;
      RECT 0 108.1 7.4 110 ;
    LAYER RDL SPACING 2 ;
      RECT 0 -20 65 -5 ;
      RECT 0 72 65 110 ;
      RECT 3 4.5 62 63.5 ;
  END
END P65_1233_PAR

MACRO P65_1233_PAR_5
  CLASS PAD ;
  ORIGIN 0 20 ;
  FOREIGN P65_1233_PAR_5 0 -20 ;
  SIZE 65 BY 130 ;
  SYMMETRY X Y R90 ;
  SITE IOSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA2 ;
    ANTENNAPARTIALCUTAREA 3.645 LAYER VIA4 ;
    PORT
      LAYER MET5 ;
        RECT 8 109 57 110 ;
      LAYER MET4 ;
        RECT 8 109 57 110 ;
      LAYER MET3 ;
        RECT 8 109 57 110 ;
      LAYER MET2 ;
        RECT 8 98.085 57 110 ;
        RECT 45.92 89.5 57 110 ;
        RECT 8 89.5 19 110 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET2 ;
        RECT 0 99.98 6.5 107.02 ;
        RECT 0 99.937 6.46 107.063 ;
        RECT 0 99.891 6.414 107.109 ;
        RECT 0 99.845 6.368 107.155 ;
        RECT 0 99.799 6.322 107.201 ;
        RECT 0 99.753 6.276 107.247 ;
        RECT 0 99.707 6.23 107.293 ;
        RECT 0 99.661 6.184 107.339 ;
        RECT 0 99.615 6.138 107.385 ;
        RECT 0 99.569 6.092 107.431 ;
        RECT 0 99.523 6.046 107.477 ;
        RECT 0 99.5 6 107.5 ;
    END
    PORT
      CLASS CORE ;
      LAYER MET5 ;
        RECT 0 99.5 65 107.5 ;
      LAYER MET4 ;
        RECT 0 99.5 65 107.5 ;
      LAYER MET3 ;
        RECT 0 99.5 65 107.5 ;
    END
  END VDD
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET5 ;
        RECT 0 68.5 65 77 ;
        RECT 0 30.788 1.5 42.212 ;
        RECT 0 30.753 1.476 42.247 ;
        RECT 0 30.707 1.43 42.293 ;
        RECT 0 30.661 1.384 42.339 ;
        RECT 0 30.615 1.338 42.385 ;
        RECT 0 30.569 1.292 42.431 ;
        RECT 0 30.523 1.246 42.477 ;
        RECT 0 30.5 1.2 42.5 ;
        RECT 0 44.288 1.5 55.712 ;
        RECT 0 44.253 1.476 55.747 ;
        RECT 0 44.207 1.43 55.793 ;
        RECT 0 44.161 1.384 55.839 ;
        RECT 0 44.115 1.338 55.885 ;
        RECT 0 44.069 1.292 55.931 ;
        RECT 0 44.023 1.246 55.977 ;
        RECT 0 44 1.2 56 ;
        RECT 0 57.788 1.5 63.212 ;
        RECT 0 57.753 1.476 63.247 ;
        RECT 0 57.707 1.43 63.293 ;
        RECT 0 57.661 1.384 63.339 ;
        RECT 0 57.615 1.338 63.385 ;
        RECT 0 57.569 1.292 63.431 ;
        RECT 0 57.523 1.246 63.477 ;
        RECT 0 57.5 1.2 63.5 ;
      LAYER MET4 ;
        RECT 0 68.5 65 77 ;
        RECT 0 30.788 1.5 42.212 ;
        RECT 0 30.753 1.476 42.247 ;
        RECT 0 30.707 1.43 42.293 ;
        RECT 0 30.661 1.384 42.339 ;
        RECT 0 30.615 1.338 42.385 ;
        RECT 0 30.569 1.292 42.431 ;
        RECT 0 30.523 1.246 42.477 ;
        RECT 0 30.5 1.2 42.5 ;
        RECT 0 44.288 1.5 55.712 ;
        RECT 0 44.253 1.476 55.747 ;
        RECT 0 44.207 1.43 55.793 ;
        RECT 0 44.161 1.384 55.839 ;
        RECT 0 44.115 1.338 55.885 ;
        RECT 0 44.069 1.292 55.931 ;
        RECT 0 44.023 1.246 55.977 ;
        RECT 0 44 1.2 56 ;
        RECT 0 57.788 1.5 63.212 ;
        RECT 0 57.753 1.476 63.247 ;
        RECT 0 57.707 1.43 63.293 ;
        RECT 0 57.661 1.384 63.339 ;
        RECT 0 57.615 1.338 63.385 ;
        RECT 0 57.569 1.292 63.431 ;
        RECT 0 57.523 1.246 63.477 ;
        RECT 0 57.5 1.2 63.5 ;
      LAYER MET3 ;
        RECT 0 68.5 65 77 ;
        RECT 0 30.788 1.5 42.212 ;
        RECT 0 30.753 1.476 42.247 ;
        RECT 0 30.707 1.43 42.293 ;
        RECT 0 30.661 1.384 42.339 ;
        RECT 0 30.615 1.338 42.385 ;
        RECT 0 30.569 1.292 42.431 ;
        RECT 0 30.523 1.246 42.477 ;
        RECT 0 30.5 1.2 42.5 ;
        RECT 0 44.288 1.5 55.712 ;
        RECT 0 44.253 1.476 55.747 ;
        RECT 0 44.207 1.43 55.793 ;
        RECT 0 44.161 1.384 55.839 ;
        RECT 0 44.115 1.338 55.885 ;
        RECT 0 44.069 1.292 55.931 ;
        RECT 0 44.023 1.246 55.977 ;
        RECT 0 44 1.2 56 ;
        RECT 0 57.788 1.5 63.212 ;
        RECT 0 57.753 1.476 63.247 ;
        RECT 0 57.707 1.43 63.293 ;
        RECT 0 57.661 1.384 63.339 ;
        RECT 0 57.615 1.338 63.385 ;
        RECT 0 57.569 1.292 63.431 ;
        RECT 0 57.523 1.246 63.477 ;
        RECT 0 57.5 1.2 63.5 ;
      LAYER MET2 ;
        RECT 0 68.5 65 77 ;
        RECT 0 57.5 65 63.5 ;
        RECT 0 44 65 56 ;
        RECT 0 30.5 65 42.5 ;
        RECT 57.015 30.5 58.205 77 ;
        RECT 51.435 30.5 52.625 77 ;
        RECT 45.855 30.5 47.045 77 ;
        RECT 40.275 30.5 41.465 77 ;
        RECT 34.695 30.5 35.885 77 ;
        RECT 29.115 30.5 30.305 77 ;
        RECT 23.535 30.5 24.725 77 ;
        RECT 17.955 30.5 19.145 77 ;
        RECT 12.375 30.5 13.565 77 ;
        RECT 6.795 30.5 7.985 77 ;
    END
  END VDDA
  PIN VSS
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 45.25 LAYER MET2 ;
    ANTENNAPARTIALCUTAREA 6.2694 LAYER VIA4 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 1.6848 LAYER VIA2 ;
    PORT
      LAYER MET5 ;
        RECT 0 91 65 98 ;
      LAYER MET4 ;
        RECT 0 91 65 98 ;
      LAYER MET3 ;
        RECT 0 91 65 98 ;
      LAYER MET2 ;
        RECT 0 91.48 6.5 97.52 ;
        RECT 0 91.437 6.46 97.563 ;
        RECT 0 91.391 6.414 97.609 ;
        RECT 0 91.345 6.368 97.655 ;
        RECT 0 91.299 6.322 97.701 ;
        RECT 0 91.253 6.276 97.747 ;
        RECT 0 91.207 6.23 97.793 ;
        RECT 0 91.161 6.184 97.839 ;
        RECT 0 91.115 6.138 97.885 ;
        RECT 0 91.069 6.092 97.931 ;
        RECT 0 91.023 6.046 97.977 ;
        RECT 0 91 6 98 ;
    END
  END VSS
  PIN VSSA
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA2 ;
    ANTENNAPARTIALCUTAREA 9.7524 LAYER VIA4 ;
    PORT
      LAYER MET5 ;
        RECT 0 78.5 65 89.5 ;
        RECT 0 3.788 1.5 15.212 ;
        RECT 0 3.753 1.476 15.247 ;
        RECT 0 3.707 1.43 15.293 ;
        RECT 0 3.661 1.384 15.339 ;
        RECT 0 3.615 1.338 15.385 ;
        RECT 0 3.569 1.292 15.431 ;
        RECT 0 3.523 1.246 15.477 ;
        RECT 0 3.5 1.2 15.5 ;
        RECT 0 17.288 1.5 28.712 ;
        RECT 0 17.253 1.476 28.747 ;
        RECT 0 17.207 1.43 28.793 ;
        RECT 0 17.161 1.384 28.839 ;
        RECT 0 17.115 1.338 28.885 ;
        RECT 0 17.069 1.292 28.931 ;
        RECT 0 17.023 1.246 28.977 ;
        RECT 0 17 1.2 29 ;
      LAYER MET4 ;
        RECT 0 78.5 65 89.5 ;
        RECT 0 3.788 1.5 15.212 ;
        RECT 0 3.753 1.476 15.247 ;
        RECT 0 3.707 1.43 15.293 ;
        RECT 0 3.661 1.384 15.339 ;
        RECT 0 3.615 1.338 15.385 ;
        RECT 0 3.569 1.292 15.431 ;
        RECT 0 3.523 1.246 15.477 ;
        RECT 0 3.5 1.2 15.5 ;
        RECT 0 17.288 1.5 28.712 ;
        RECT 0 17.253 1.476 28.747 ;
        RECT 0 17.207 1.43 28.793 ;
        RECT 0 17.161 1.384 28.839 ;
        RECT 0 17.115 1.338 28.885 ;
        RECT 0 17.069 1.292 28.931 ;
        RECT 0 17.023 1.246 28.977 ;
        RECT 0 17 1.2 29 ;
      LAYER MET3 ;
        RECT 0 78.5 65 89.5 ;
        RECT 0 3.788 1.5 15.212 ;
        RECT 0 3.753 1.476 15.247 ;
        RECT 0 3.707 1.43 15.293 ;
        RECT 0 3.661 1.384 15.339 ;
        RECT 0 3.615 1.338 15.385 ;
        RECT 0 3.569 1.292 15.431 ;
        RECT 0 3.523 1.246 15.477 ;
        RECT 0 3.5 1.2 15.5 ;
        RECT 0 17.288 1.5 28.712 ;
        RECT 0 17.253 1.476 28.747 ;
        RECT 0 17.207 1.43 28.793 ;
        RECT 0 17.161 1.384 28.839 ;
        RECT 0 17.115 1.338 28.885 ;
        RECT 0 17.069 1.292 28.931 ;
        RECT 0 17.023 1.246 28.977 ;
        RECT 0 17 1.2 29 ;
      LAYER MET2 ;
        RECT 0 17 65 29 ;
        RECT 0 3.5 65 15.5 ;
        RECT 59.805 3.5 60.995 29 ;
        RECT 54.225 3.5 55.415 29 ;
        RECT 48.645 3.5 49.835 29 ;
        RECT 43.065 3.5 44.255 29 ;
        RECT 37.485 3.5 38.675 29 ;
        RECT 31.905 3.5 33.095 29 ;
        RECT 26.325 3.5 27.515 29 ;
        RECT 20.745 3.5 21.935 29 ;
        RECT 15.165 3.5 16.355 29 ;
        RECT 9.585 3.5 10.775 29 ;
        RECT 4.005 3.5 5.195 29 ;
        RECT 0 78.98 6.5 89.02 ;
        RECT 0 78.937 6.46 89.063 ;
        RECT 0 78.891 6.414 89.109 ;
        RECT 0 78.845 6.368 89.155 ;
        RECT 0 78.799 6.322 89.201 ;
        RECT 0 78.753 6.276 89.247 ;
        RECT 0 78.707 6.23 89.293 ;
        RECT 0 78.661 6.184 89.339 ;
        RECT 0 78.615 6.138 89.385 ;
        RECT 0 78.569 6.092 89.431 ;
        RECT 0 78.523 6.046 89.477 ;
        RECT 0 78.5 6 89.5 ;
    END
  END VSSA
  PIN PAD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER T4M2 ;
        RECT 57 0.983 62 66.017 ;
        RECT 57 0.943 61.966 66.057 ;
        RECT 57 0.897 61.92 66.103 ;
        RECT 57 0.851 61.874 66.149 ;
        RECT 57 0.805 61.828 66.195 ;
        RECT 57 0.759 61.782 66.241 ;
        RECT 57 0.713 61.736 66.287 ;
        RECT 57 0.667 61.69 66.333 ;
        RECT 57 0.621 61.644 66.379 ;
        RECT 57 0.575 61.598 66.425 ;
        RECT 57 0.529 61.552 66.471 ;
        RECT 57 0.483 61.506 66.517 ;
        RECT 57 0.437 61.46 66.563 ;
        RECT 57 0.391 61.414 66.609 ;
        RECT 57 0.345 61.368 66.655 ;
        RECT 57 0.299 61.322 66.701 ;
        RECT 57 0.253 61.276 66.747 ;
        RECT 57 0.207 61.23 66.793 ;
        RECT 57 0.161 61.184 66.839 ;
        RECT 57 0.115 61.138 66.885 ;
        RECT 57 0.069 61.092 66.931 ;
        RECT 57 0.023 61.046 66.977 ;
        RECT 4 57.5 61 67 ;
        RECT 3 43.5 62 51 ;
        RECT 3 29.5 62 37 ;
        RECT 3 15.5 62 23 ;
        RECT 4 0 61 9 ;
        RECT 43 0 50.5 67 ;
        RECT 29 0 36.5 67 ;
        RECT 15 0 22.5 67 ;
        RECT 3 0.977 8.5 66.023 ;
        RECT 3.966 0.017 8.5 66.983 ;
        RECT 3.92 0.057 8.5 66.943 ;
        RECT 3.874 0.103 8.5 66.897 ;
        RECT 3.828 0.149 8.5 66.851 ;
        RECT 3.782 0.195 8.5 66.805 ;
        RECT 3.736 0.241 8.5 66.759 ;
        RECT 3.69 0.287 8.5 66.713 ;
        RECT 3.644 0.333 8.5 66.667 ;
        RECT 3.598 0.379 8.5 66.621 ;
        RECT 3.552 0.425 8.5 66.575 ;
        RECT 3.506 0.471 8.5 66.529 ;
        RECT 3.46 0.517 8.5 66.483 ;
        RECT 3.414 0.563 8.5 66.437 ;
        RECT 3.368 0.609 8.5 66.391 ;
        RECT 3.322 0.655 8.5 66.345 ;
        RECT 3.276 0.701 8.5 66.299 ;
        RECT 3.23 0.747 8.5 66.253 ;
        RECT 3.184 0.793 8.5 66.207 ;
        RECT 3.138 0.839 8.5 66.161 ;
        RECT 3.092 0.885 8.5 66.115 ;
        RECT 3.046 0.931 8.5 66.069 ;
    END
  END PAD
  OBS
    LAYER MET1 SPACING 0.09 ;
      RECT 0 -20 65 110 ;
    LAYER MET2 SPACING 0.1 ;
      RECT 57.175 77.175 65 110 ;
      RECT 0 107.675 7.825 110 ;
      RECT 6.675 77.175 7.825 110 ;
      RECT 6.175 107.652 7.825 110 ;
      RECT 6.635 107.195 7.825 110 ;
      RECT 6.221 107.606 7.825 110 ;
      RECT 6.589 107.238 7.825 110 ;
      RECT 6.267 107.56 7.825 110 ;
      RECT 6.543 107.284 7.825 110 ;
      RECT 6.313 107.514 7.825 110 ;
      RECT 6.497 107.33 7.825 110 ;
      RECT 6.359 107.468 7.825 110 ;
      RECT 6.451 107.376 7.825 110 ;
      RECT 6.405 107.422 7.825 110 ;
      RECT 6.635 97.695 7.825 99.805 ;
      RECT 6.589 97.738 7.825 99.762 ;
      RECT 6.543 97.784 7.825 99.716 ;
      RECT 6.497 97.83 7.825 99.67 ;
      RECT 6.451 97.876 7.825 99.624 ;
      RECT 6.405 97.922 7.825 99.578 ;
      RECT 6.359 97.968 7.825 99.532 ;
      RECT 6.313 98.014 7.825 99.486 ;
      RECT 6.267 98.06 7.825 99.44 ;
      RECT 6.221 98.106 7.825 99.394 ;
      RECT 6.175 98.152 7.825 99.348 ;
      RECT 0 98.175 7.825 99.325 ;
      RECT 19.175 77.175 45.745 97.91 ;
      RECT 6.635 89.195 7.825 91.305 ;
      RECT 6.589 89.238 7.825 91.262 ;
      RECT 6.543 89.284 7.825 91.216 ;
      RECT 6.497 89.33 7.825 91.17 ;
      RECT 6.451 89.376 7.825 91.124 ;
      RECT 6.405 89.422 7.825 91.078 ;
      RECT 6.359 89.468 7.825 91.032 ;
      RECT 6.313 89.514 7.825 90.986 ;
      RECT 6.267 89.56 7.825 90.94 ;
      RECT 6.221 89.606 7.825 90.894 ;
      RECT 6.175 89.652 7.825 90.848 ;
      RECT 0 89.675 7.825 90.825 ;
      RECT 6.675 77.175 65 89.325 ;
      RECT 6.635 77.175 65 78.805 ;
      RECT 6.589 77.175 65 78.762 ;
      RECT 6.543 77.175 65 78.716 ;
      RECT 6.497 77.175 65 78.67 ;
      RECT 6.451 77.175 65 78.624 ;
      RECT 6.405 77.175 65 78.578 ;
      RECT 6.359 77.175 65 78.532 ;
      RECT 6.313 77.175 65 78.486 ;
      RECT 6.267 77.175 65 78.44 ;
      RECT 6.221 77.175 65 78.394 ;
      RECT 6.175 77.175 65 78.348 ;
      RECT 0 77.175 65 78.325 ;
      RECT 0 -20 65 3.325 ;
      RECT 61.17 15.675 65 16.825 ;
      RECT 0 29.175 65 30.325 ;
      RECT 58.38 42.675 65 43.825 ;
      RECT 58.38 56.175 65 57.325 ;
      RECT 58.38 63.675 65 68.325 ;
      RECT 55.59 15.675 59.63 16.825 ;
      RECT 52.8 42.675 56.84 43.825 ;
      RECT 52.8 56.175 56.84 57.325 ;
      RECT 52.8 63.675 56.84 68.325 ;
      RECT 50.01 15.675 54.05 16.825 ;
      RECT 47.22 42.675 51.26 43.825 ;
      RECT 47.22 56.175 51.26 57.325 ;
      RECT 47.22 63.675 51.26 68.325 ;
      RECT 44.43 15.675 48.47 16.825 ;
      RECT 41.64 42.675 45.68 43.825 ;
      RECT 41.64 56.175 45.68 57.325 ;
      RECT 41.64 63.675 45.68 68.325 ;
      RECT 38.85 15.675 42.89 16.825 ;
      RECT 36.06 42.675 40.1 43.825 ;
      RECT 36.06 56.175 40.1 57.325 ;
      RECT 36.06 63.675 40.1 68.325 ;
      RECT 33.27 15.675 37.31 16.825 ;
      RECT 30.48 42.675 34.52 43.825 ;
      RECT 30.48 56.175 34.52 57.325 ;
      RECT 30.48 63.675 34.52 68.325 ;
      RECT 27.69 15.675 31.73 16.825 ;
      RECT 24.9 42.675 28.94 43.825 ;
      RECT 24.9 56.175 28.94 57.325 ;
      RECT 24.9 63.675 28.94 68.325 ;
      RECT 22.11 15.675 26.15 16.825 ;
      RECT 19.32 42.675 23.36 43.825 ;
      RECT 19.32 56.175 23.36 57.325 ;
      RECT 19.32 63.675 23.36 68.325 ;
      RECT 16.53 15.675 20.57 16.825 ;
      RECT 13.74 42.675 17.78 43.825 ;
      RECT 13.74 56.175 17.78 57.325 ;
      RECT 13.74 63.675 17.78 68.325 ;
      RECT 10.95 15.675 14.99 16.825 ;
      RECT 8.16 42.675 12.2 43.825 ;
      RECT 8.16 56.175 12.2 57.325 ;
      RECT 8.16 63.675 12.2 68.325 ;
      RECT 5.37 15.675 9.41 16.825 ;
      RECT 0 42.675 6.62 43.825 ;
      RECT 0 56.175 6.62 57.325 ;
      RECT 0 63.675 6.62 68.325 ;
      RECT 0 15.675 3.83 16.825 ;
    LAYER MET3 SPACING 0.1 ;
      RECT 58.37 63.665 65 68.325 ;
      RECT 52.79 57.5 56.85 68.325 ;
      RECT 47.21 57.5 51.27 68.325 ;
      RECT 41.63 57.5 45.69 68.325 ;
      RECT 36.05 57.5 40.11 68.325 ;
      RECT 30.47 -20 34.53 68.325 ;
      RECT 24.89 57.5 28.95 68.325 ;
      RECT 19.31 57.5 23.37 68.325 ;
      RECT 13.73 57.5 17.79 68.325 ;
      RECT 8.15 57.5 12.21 68.325 ;
      RECT 0 63.675 6.63 68.325 ;
      RECT 57 -20 62 67 ;
      RECT 1.375 63.665 65 67 ;
      RECT 3 57.5 62 67 ;
      RECT 43 -20 50.5 67 ;
      RECT 29 -20 36.5 67 ;
      RECT 15 -20 22.5 67 ;
      RECT 3 -20 8.5 67 ;
      RECT 57 56.165 65 57.335 ;
      RECT 41.63 56.165 51.27 57.335 ;
      RECT 24.89 56.165 40.11 57.335 ;
      RECT 13.73 56.165 23.37 57.335 ;
      RECT 1.375 56.165 12.21 57.335 ;
      RECT 0 56.175 12.21 57.325 ;
      RECT 3 43.5 62 51 ;
      RECT 57 42.665 65 43.835 ;
      RECT 0 42.675 12.21 43.825 ;
      RECT 52.79 42.665 56.85 51 ;
      RECT 41.63 42.665 51.27 51 ;
      RECT 24.89 42.665 40.11 51 ;
      RECT 13.73 42.665 23.37 51 ;
      RECT 1.375 42.665 12.21 43.835 ;
      RECT 3 29.165 62 37 ;
      RECT 1.375 29.165 65 30.335 ;
      RECT 0 29.175 65 30.325 ;
      RECT 3 15.5 62 23 ;
      RECT 1.375 15.665 65 16.835 ;
      RECT 0 15.675 65 16.825 ;
      RECT 3 -20 62 9 ;
      RECT 1.375 -20 65 3.335 ;
      RECT 0 -20 65 3.325 ;
      RECT 63.8 3.5 65 15.5 ;
      RECT 63.776 3.512 65 15.488 ;
      RECT 63.73 3.547 65 15.453 ;
      RECT 63.684 3.593 65 15.407 ;
      RECT 63.638 3.639 65 15.361 ;
      RECT 63.592 3.685 65 15.315 ;
      RECT 63.546 3.731 65 15.269 ;
      RECT 63.5 3.777 65 15.223 ;
      RECT 63.8 17 65 29 ;
      RECT 63.776 17.012 65 28.988 ;
      RECT 63.73 17.047 65 28.953 ;
      RECT 63.684 17.093 65 28.907 ;
      RECT 63.638 17.139 65 28.861 ;
      RECT 63.592 17.185 65 28.815 ;
      RECT 63.546 17.231 65 28.769 ;
      RECT 63.5 17.277 65 28.723 ;
      RECT 63.8 30.5 65 42.5 ;
      RECT 63.776 30.512 65 42.488 ;
      RECT 63.73 30.547 65 42.453 ;
      RECT 63.684 30.593 65 42.407 ;
      RECT 63.638 30.639 65 42.361 ;
      RECT 63.592 30.685 65 42.315 ;
      RECT 63.546 30.731 65 42.269 ;
      RECT 63.5 30.777 65 42.223 ;
      RECT 63.8 44 65 56 ;
      RECT 63.776 44.012 65 55.988 ;
      RECT 63.73 44.047 65 55.953 ;
      RECT 63.684 44.093 65 55.907 ;
      RECT 63.638 44.139 65 55.861 ;
      RECT 63.592 44.185 65 55.815 ;
      RECT 63.546 44.231 65 55.769 ;
      RECT 63.5 44.277 65 55.723 ;
      RECT 63.8 57.5 65 63.5 ;
      RECT 63.776 57.512 65 63.488 ;
      RECT 63.73 57.547 65 63.453 ;
      RECT 63.684 57.593 65 63.407 ;
      RECT 63.638 57.639 65 63.361 ;
      RECT 63.592 57.685 65 63.315 ;
      RECT 63.546 57.731 65 63.269 ;
      RECT 63.5 57.777 65 63.223 ;
      RECT 57.175 107.675 65 110 ;
      RECT 57.165 107.675 65 108.825 ;
      RECT 0 107.675 7.825 110 ;
      RECT 0 107.675 7.835 108.825 ;
      RECT 0 77.175 65 78.325 ;
      RECT 57.165 89.675 65 90.825 ;
      RECT 57.165 98.175 65 99.325 ;
      RECT 52.79 56.165 56.85 57.335 ;
      RECT 19.165 89.675 45.755 90.825 ;
      RECT 0 89.675 7.835 90.825 ;
      RECT 0 98.175 7.835 99.325 ;
    LAYER MET4 SPACING 0.1 ;
      RECT 0 63.675 65 68.325 ;
      RECT 1.675 -20 65 68.325 ;
      RECT 1.375 63.652 65 68.325 ;
      RECT 1.651 63.387 65 68.325 ;
      RECT 1.421 63.606 65 68.325 ;
      RECT 1.605 63.422 65 68.325 ;
      RECT 1.467 63.56 65 68.325 ;
      RECT 1.559 63.468 65 68.325 ;
      RECT 1.513 63.514 65 68.325 ;
      RECT 1.651 55.887 65 57.613 ;
      RECT 1.605 55.922 65 57.578 ;
      RECT 1.559 55.968 65 57.532 ;
      RECT 1.513 56.014 65 57.486 ;
      RECT 1.467 56.06 65 57.44 ;
      RECT 1.421 56.106 65 57.394 ;
      RECT 1.375 56.152 65 57.348 ;
      RECT 0 56.175 65 57.325 ;
      RECT 1.651 42.387 65 44.113 ;
      RECT 1.605 42.422 65 44.078 ;
      RECT 1.559 42.468 65 44.032 ;
      RECT 1.513 42.514 65 43.986 ;
      RECT 1.467 42.56 65 43.94 ;
      RECT 1.421 42.606 65 43.894 ;
      RECT 1.375 42.652 65 43.848 ;
      RECT 0 42.675 65 43.825 ;
      RECT 1.651 28.887 65 30.613 ;
      RECT 1.605 28.922 65 30.578 ;
      RECT 1.559 28.968 65 30.532 ;
      RECT 1.513 29.014 65 30.486 ;
      RECT 1.467 29.06 65 30.44 ;
      RECT 1.421 29.106 65 30.394 ;
      RECT 1.375 29.152 65 30.348 ;
      RECT 0 29.175 65 30.325 ;
      RECT 1.651 15.387 65 17.113 ;
      RECT 1.605 15.422 65 17.078 ;
      RECT 1.559 15.468 65 17.032 ;
      RECT 1.513 15.514 65 16.986 ;
      RECT 1.467 15.56 65 16.94 ;
      RECT 1.421 15.606 65 16.894 ;
      RECT 1.375 15.652 65 16.848 ;
      RECT 0 15.675 65 16.825 ;
      RECT 1.651 -20 65 3.613 ;
      RECT 1.605 -20 65 3.578 ;
      RECT 1.559 -20 65 3.532 ;
      RECT 1.513 -20 65 3.486 ;
      RECT 1.467 -20 65 3.44 ;
      RECT 1.421 -20 65 3.394 ;
      RECT 1.375 -20 65 3.348 ;
      RECT 0 -20 65 3.325 ;
      RECT 57.175 107.675 65 110 ;
      RECT 0 107.675 7.825 110 ;
      RECT 0 107.675 65 108.825 ;
      RECT 0 77.175 65 78.325 ;
      RECT 0 89.675 65 90.825 ;
      RECT 0 98.175 65 99.325 ;
    LAYER MET5 SPACING 0.1 ;
      RECT 0 63.83 65 68.17 ;
      RECT 1.83 -20 65 68.17 ;
      RECT 1.53 63.807 65 68.17 ;
      RECT 1.806 63.542 65 68.17 ;
      RECT 1.576 63.761 65 68.17 ;
      RECT 1.76 63.577 65 68.17 ;
      RECT 1.622 63.715 65 68.17 ;
      RECT 1.714 63.623 65 68.17 ;
      RECT 1.668 63.669 65 68.17 ;
      RECT 1.806 56.042 65 57.458 ;
      RECT 1.76 56.077 65 57.423 ;
      RECT 1.714 56.123 65 57.377 ;
      RECT 1.668 56.169 65 57.331 ;
      RECT 1.622 56.215 65 57.285 ;
      RECT 1.576 56.261 65 57.239 ;
      RECT 1.53 56.307 65 57.193 ;
      RECT 0 56.33 65 57.17 ;
      RECT 1.806 42.542 65 43.958 ;
      RECT 1.76 42.577 65 43.923 ;
      RECT 1.714 42.623 65 43.877 ;
      RECT 1.668 42.669 65 43.831 ;
      RECT 1.622 42.715 65 43.785 ;
      RECT 1.576 42.761 65 43.739 ;
      RECT 1.53 42.807 65 43.693 ;
      RECT 0 42.83 65 43.67 ;
      RECT 1.806 29.042 65 30.458 ;
      RECT 1.76 29.077 65 30.423 ;
      RECT 1.714 29.123 65 30.377 ;
      RECT 1.668 29.169 65 30.331 ;
      RECT 1.622 29.215 65 30.285 ;
      RECT 1.576 29.261 65 30.239 ;
      RECT 1.53 29.307 65 30.193 ;
      RECT 0 29.33 65 30.17 ;
      RECT 1.806 15.542 65 16.958 ;
      RECT 1.76 15.577 65 16.923 ;
      RECT 1.714 15.623 65 16.877 ;
      RECT 1.668 15.669 65 16.831 ;
      RECT 1.622 15.715 65 16.785 ;
      RECT 1.576 15.761 65 16.739 ;
      RECT 1.53 15.807 65 16.693 ;
      RECT 0 15.83 65 16.67 ;
      RECT 1.806 -20 65 3.458 ;
      RECT 1.76 -20 65 3.423 ;
      RECT 1.714 -20 65 3.377 ;
      RECT 1.668 -20 65 3.331 ;
      RECT 1.622 -20 65 3.285 ;
      RECT 1.576 -20 65 3.239 ;
      RECT 1.53 -20 65 3.193 ;
      RECT 0 -20 65 3.17 ;
      RECT 57.33 107.83 65 110 ;
      RECT 0 107.83 7.67 110 ;
      RECT 0 107.83 65 108.67 ;
      RECT 0 77.33 65 78.17 ;
      RECT 0 89.83 65 90.67 ;
      RECT 0 98.33 65 99.17 ;
    LAYER T4M2 SPACING 0.4 ;
      RECT 64.584 -20 65 -3.193 ;
      RECT 0 -20 0.428 -3.205 ;
      RECT 64.538 -20 65 -3.239 ;
      RECT 0 -20 0.474 -3.251 ;
      RECT 64.492 -20 65 -3.285 ;
      RECT 0 -20 0.52 -3.297 ;
      RECT 64.446 -20 65 -3.331 ;
      RECT 0 -20 0.566 -3.343 ;
      RECT 64.4 -20 65 -3.377 ;
      RECT 0 -20 0.6 -3.383 ;
      RECT 0 -20 65 -3.4 ;
      RECT 57.6 108.1 65 110 ;
      RECT 0 108.1 7.4 110 ;
    LAYER RDL SPACING 2 ;
      RECT 0 -20 65 -5 ;
      RECT 0 72 65 110 ;
      RECT 3 4.5 62 63.5 ;
  END
END P65_1233_PAR_5

MACRO P65_1233_PBMUX
  CLASS PAD ;
  ORIGIN 0 20 ;
  FOREIGN P65_1233_PBMUX 0 -20 ;
  SIZE 65 BY 130 ;
  SYMMETRY X Y R90 ;
  SITE IOSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA2 ;
    ANTENNAPARTIALCUTAREA 0.0486 LAYER VIA4 ;
    PORT
      LAYER MET5 ;
        RECT 60.64 109.4 61.84 110 ;
      LAYER MET4 ;
        RECT 60.64 109.4 61.84 110 ;
      LAYER MET3 ;
        RECT 60.64 109.4 61.84 110 ;
      LAYER MET2 ;
        RECT 60.64 109.4 61.84 110 ;
    END
  END A
  PIN C
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA2 ;
    ANTENNAPARTIALCUTAREA 0.0486 LAYER VIA4 ;
    PORT
      LAYER MET5 ;
        RECT 44.31 109.4 45.51 110 ;
      LAYER MET4 ;
        RECT 44.31 109.4 45.51 110 ;
      LAYER MET3 ;
        RECT 44.31 109.4 45.51 110 ;
      LAYER MET2 ;
        RECT 44.31 109.4 45.51 110 ;
    END
  END C
  PIN CS
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA2 ;
    ANTENNAPARTIALCUTAREA 0.0486 LAYER VIA4 ;
    PORT
      LAYER MET5 ;
        RECT 28.87 109.4 30.07 110 ;
      LAYER MET4 ;
        RECT 28.87 109.4 30.07 110 ;
      LAYER MET3 ;
        RECT 28.87 109.4 30.07 110 ;
      LAYER MET2 ;
        RECT 28.87 109.4 30.07 110 ;
    END
  END CS
  PIN DS0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA2 ;
    ANTENNAPARTIALCUTAREA 0.0486 LAYER VIA4 ;
    PORT
      LAYER MET5 ;
        RECT 8.325 109.4 9.525 110 ;
      LAYER MET4 ;
        RECT 8.325 109.4 9.525 110 ;
      LAYER MET3 ;
        RECT 8.325 109.4 9.525 110 ;
      LAYER MET2 ;
        RECT 8.325 109.4 9.525 110 ;
    END
  END DS0
  PIN DS1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA2 ;
    ANTENNAPARTIALCUTAREA 0.0486 LAYER VIA4 ;
    PORT
      LAYER MET5 ;
        RECT 14.185 109.4 15.385 110 ;
      LAYER MET4 ;
        RECT 14.185 109.4 15.385 110 ;
      LAYER MET3 ;
        RECT 14.185 109.4 15.385 110 ;
      LAYER MET2 ;
        RECT 14.185 109.4 15.385 110 ;
    END
  END DS1
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA2 ;
    ANTENNAPARTIALCUTAREA 0.0486 LAYER VIA4 ;
    PORT
      LAYER MET5 ;
        RECT 49.455 109.4 50.655 110 ;
      LAYER MET4 ;
        RECT 49.455 109.4 50.655 110 ;
      LAYER MET3 ;
        RECT 49.455 109.4 50.655 110 ;
      LAYER MET2 ;
        RECT 49.455 109.4 50.655 110 ;
    END
  END I
  PIN IE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8141 LAYER MET2 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA2 ;
    ANTENNAPARTIALCUTAREA 0.0486 LAYER VIA4 ;
    PORT
      LAYER MET5 ;
        RECT 37.035 109.4 38.235 110 ;
      LAYER MET4 ;
        RECT 37.035 109.4 38.235 110 ;
      LAYER MET3 ;
        RECT 37.035 109.4 38.235 110 ;
      LAYER MET2 ;
        RECT 37.035 109.4 38.235 110 ;
    END
  END IE
  PIN OD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5411 LAYER MET2 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA2 ;
    ANTENNAPARTIALCUTAREA 0.0486 LAYER VIA4 ;
    PORT
      LAYER MET5 ;
        RECT 5.65 109.4 6.85 110 ;
      LAYER MET4 ;
        RECT 5.65 109.4 6.85 110 ;
      LAYER MET3 ;
        RECT 5.65 109.4 6.85 110 ;
      LAYER MET2 ;
        RECT 5.65 109.4 6.85 110 ;
    END
  END OD
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA2 ;
    ANTENNAPARTIALCUTAREA 0.0486 LAYER VIA4 ;
    PORT
      LAYER MET5 ;
        RECT 46.87 109.4 48.07 110 ;
      LAYER MET4 ;
        RECT 46.87 109.4 48.07 110 ;
      LAYER MET3 ;
        RECT 46.87 109.4 48.07 110 ;
      LAYER MET2 ;
        RECT 46.87 109.4 48.07 110 ;
    END
  END OE
  PIN PD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA2 ;
    ANTENNAPARTIALCUTAREA 0.0486 LAYER VIA4 ;
    PORT
      LAYER MET5 ;
        RECT 25.94 109.4 27.14 110 ;
      LAYER MET4 ;
        RECT 25.94 109.4 27.14 110 ;
      LAYER MET3 ;
        RECT 25.94 109.4 27.14 110 ;
      LAYER MET2 ;
        RECT 25.94 109.4 27.14 110 ;
    END
  END PD
  PIN PU
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA2 ;
    ANTENNAPARTIALCUTAREA 0.0486 LAYER VIA4 ;
    PORT
      LAYER MET5 ;
        RECT 21.395 109.4 22.595 110 ;
      LAYER MET4 ;
        RECT 21.395 109.4 22.595 110 ;
      LAYER MET3 ;
        RECT 21.395 109.4 22.595 110 ;
      LAYER MET2 ;
        RECT 21.395 109.4 22.595 110 ;
    END
  END PU
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER MET5 ;
        RECT 0 99.5 65 107.5 ;
      LAYER MET4 ;
        RECT 0 99.5 65 107.5 ;
      LAYER MET3 ;
        RECT 0 99.5 65 107.5 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET5 ;
        RECT 0 68.5 65 77 ;
        RECT 0 30.788 1.5 42.212 ;
        RECT 0 30.753 1.476 42.247 ;
        RECT 0 30.707 1.43 42.293 ;
        RECT 0 30.661 1.384 42.339 ;
        RECT 0 30.615 1.338 42.385 ;
        RECT 0 30.569 1.292 42.431 ;
        RECT 0 30.523 1.246 42.477 ;
        RECT 0 30.5 1.2 42.5 ;
        RECT 0 44.288 1.5 55.712 ;
        RECT 0 44.253 1.476 55.747 ;
        RECT 0 44.207 1.43 55.793 ;
        RECT 0 44.161 1.384 55.839 ;
        RECT 0 44.115 1.338 55.885 ;
        RECT 0 44.069 1.292 55.931 ;
        RECT 0 44.023 1.246 55.977 ;
        RECT 0 44 1.2 56 ;
        RECT 0 57.788 1.5 63.212 ;
        RECT 0 57.753 1.476 63.247 ;
        RECT 0 57.707 1.43 63.293 ;
        RECT 0 57.661 1.384 63.339 ;
        RECT 0 57.615 1.338 63.385 ;
        RECT 0 57.569 1.292 63.431 ;
        RECT 0 57.523 1.246 63.477 ;
        RECT 0 57.5 1.2 63.5 ;
      LAYER MET4 ;
        RECT 0 68.5 65 77 ;
        RECT 0 30.788 1.5 42.212 ;
        RECT 0 30.753 1.476 42.247 ;
        RECT 0 30.707 1.43 42.293 ;
        RECT 0 30.661 1.384 42.339 ;
        RECT 0 30.615 1.338 42.385 ;
        RECT 0 30.569 1.292 42.431 ;
        RECT 0 30.523 1.246 42.477 ;
        RECT 0 30.5 1.2 42.5 ;
        RECT 0 44.288 1.5 55.712 ;
        RECT 0 44.253 1.476 55.747 ;
        RECT 0 44.207 1.43 55.793 ;
        RECT 0 44.161 1.384 55.839 ;
        RECT 0 44.115 1.338 55.885 ;
        RECT 0 44.069 1.292 55.931 ;
        RECT 0 44.023 1.246 55.977 ;
        RECT 0 44 1.2 56 ;
        RECT 0 57.788 1.5 63.212 ;
        RECT 0 57.753 1.476 63.247 ;
        RECT 0 57.707 1.43 63.293 ;
        RECT 0 57.661 1.384 63.339 ;
        RECT 0 57.615 1.338 63.385 ;
        RECT 0 57.569 1.292 63.431 ;
        RECT 0 57.523 1.246 63.477 ;
        RECT 0 57.5 1.2 63.5 ;
      LAYER MET3 ;
        RECT 0 68.5 65 77 ;
        RECT 0 30.788 1.5 42.212 ;
        RECT 0 30.753 1.476 42.247 ;
        RECT 0 30.707 1.43 42.293 ;
        RECT 0 30.661 1.384 42.339 ;
        RECT 0 30.615 1.338 42.385 ;
        RECT 0 30.569 1.292 42.431 ;
        RECT 0 30.523 1.246 42.477 ;
        RECT 0 30.5 1.2 42.5 ;
        RECT 0 44.288 1.5 55.712 ;
        RECT 0 44.253 1.476 55.747 ;
        RECT 0 44.207 1.43 55.793 ;
        RECT 0 44.161 1.384 55.839 ;
        RECT 0 44.115 1.338 55.885 ;
        RECT 0 44.069 1.292 55.931 ;
        RECT 0 44.023 1.246 55.977 ;
        RECT 0 44 1.2 56 ;
        RECT 0 57.788 1.5 63.212 ;
        RECT 0 57.753 1.476 63.247 ;
        RECT 0 57.707 1.43 63.293 ;
        RECT 0 57.661 1.384 63.339 ;
        RECT 0 57.615 1.338 63.385 ;
        RECT 0 57.569 1.292 63.431 ;
        RECT 0 57.523 1.246 63.477 ;
        RECT 0 57.5 1.2 63.5 ;
    END
  END VDDIO
  PIN VSS
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 10.692 LAYER VIA4 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    PORT
      LAYER MET5 ;
        RECT 0 91 65 98 ;
      LAYER MET4 ;
        RECT 0 91 65 98 ;
      LAYER MET3 ;
        RECT 0 91 65 98 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 17.82 LAYER VIA4 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    PORT
      LAYER MET5 ;
        RECT 0 78.5 65 89.5 ;
        RECT 0 3.788 1.5 15.212 ;
        RECT 0 3.753 1.476 15.247 ;
        RECT 0 3.707 1.43 15.293 ;
        RECT 0 3.661 1.384 15.339 ;
        RECT 0 3.615 1.338 15.385 ;
        RECT 0 3.569 1.292 15.431 ;
        RECT 0 3.523 1.246 15.477 ;
        RECT 0 3.5 1.2 15.5 ;
        RECT 0 17.288 1.5 28.712 ;
        RECT 0 17.253 1.476 28.747 ;
        RECT 0 17.207 1.43 28.793 ;
        RECT 0 17.161 1.384 28.839 ;
        RECT 0 17.115 1.338 28.885 ;
        RECT 0 17.069 1.292 28.931 ;
        RECT 0 17.023 1.246 28.977 ;
        RECT 0 17 1.2 29 ;
      LAYER MET4 ;
        RECT 0 78.5 65 89.5 ;
        RECT 0 3.788 1.5 15.212 ;
        RECT 0 3.753 1.476 15.247 ;
        RECT 0 3.707 1.43 15.293 ;
        RECT 0 3.661 1.384 15.339 ;
        RECT 0 3.615 1.338 15.385 ;
        RECT 0 3.569 1.292 15.431 ;
        RECT 0 3.523 1.246 15.477 ;
        RECT 0 3.5 1.2 15.5 ;
        RECT 0 17.288 1.5 28.712 ;
        RECT 0 17.253 1.476 28.747 ;
        RECT 0 17.207 1.43 28.793 ;
        RECT 0 17.161 1.384 28.839 ;
        RECT 0 17.115 1.338 28.885 ;
        RECT 0 17.069 1.292 28.931 ;
        RECT 0 17.023 1.246 28.977 ;
        RECT 0 17 1.2 29 ;
      LAYER MET3 ;
        RECT 0 78.5 65 89.5 ;
        RECT 0 3.788 1.5 15.212 ;
        RECT 0 3.753 1.476 15.247 ;
        RECT 0 3.707 1.43 15.293 ;
        RECT 0 3.661 1.384 15.339 ;
        RECT 0 3.615 1.338 15.385 ;
        RECT 0 3.569 1.292 15.431 ;
        RECT 0 3.523 1.246 15.477 ;
        RECT 0 3.5 1.2 15.5 ;
        RECT 0 17.288 1.5 28.712 ;
        RECT 0 17.253 1.476 28.747 ;
        RECT 0 17.207 1.43 28.793 ;
        RECT 0 17.161 1.384 28.839 ;
        RECT 0 17.115 1.338 28.885 ;
        RECT 0 17.069 1.292 28.931 ;
        RECT 0 17.023 1.246 28.977 ;
        RECT 0 17 1.2 29 ;
    END
  END VSSIO
  PIN PAD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER T4M2 ;
        RECT 57 0.983 62 66.017 ;
        RECT 57 0.943 61.966 66.057 ;
        RECT 57 0.897 61.92 66.103 ;
        RECT 57 0.851 61.874 66.149 ;
        RECT 57 0.805 61.828 66.195 ;
        RECT 57 0.759 61.782 66.241 ;
        RECT 57 0.713 61.736 66.287 ;
        RECT 57 0.667 61.69 66.333 ;
        RECT 57 0.621 61.644 66.379 ;
        RECT 57 0.575 61.598 66.425 ;
        RECT 57 0.529 61.552 66.471 ;
        RECT 57 0.483 61.506 66.517 ;
        RECT 57 0.437 61.46 66.563 ;
        RECT 57 0.391 61.414 66.609 ;
        RECT 57 0.345 61.368 66.655 ;
        RECT 57 0.299 61.322 66.701 ;
        RECT 57 0.253 61.276 66.747 ;
        RECT 57 0.207 61.23 66.793 ;
        RECT 57 0.161 61.184 66.839 ;
        RECT 57 0.115 61.138 66.885 ;
        RECT 57 0.069 61.092 66.931 ;
        RECT 57 0.023 61.046 66.977 ;
        RECT 4 57.5 61 67 ;
        RECT 3 43.5 62 51 ;
        RECT 3 29.5 62 37 ;
        RECT 3 15.5 62 23 ;
        RECT 4 0 61 9 ;
        RECT 43 0 50.5 67 ;
        RECT 29 0 36.5 67 ;
        RECT 15 0 22.5 67 ;
        RECT 3 0.977 8.5 66.023 ;
        RECT 3.966 0.017 8.5 66.983 ;
        RECT 3.92 0.057 8.5 66.943 ;
        RECT 3.874 0.103 8.5 66.897 ;
        RECT 3.828 0.149 8.5 66.851 ;
        RECT 3.782 0.195 8.5 66.805 ;
        RECT 3.736 0.241 8.5 66.759 ;
        RECT 3.69 0.287 8.5 66.713 ;
        RECT 3.644 0.333 8.5 66.667 ;
        RECT 3.598 0.379 8.5 66.621 ;
        RECT 3.552 0.425 8.5 66.575 ;
        RECT 3.506 0.471 8.5 66.529 ;
        RECT 3.46 0.517 8.5 66.483 ;
        RECT 3.414 0.563 8.5 66.437 ;
        RECT 3.368 0.609 8.5 66.391 ;
        RECT 3.322 0.655 8.5 66.345 ;
        RECT 3.276 0.701 8.5 66.299 ;
        RECT 3.23 0.747 8.5 66.253 ;
        RECT 3.184 0.793 8.5 66.207 ;
        RECT 3.138 0.839 8.5 66.161 ;
        RECT 3.092 0.885 8.5 66.115 ;
        RECT 3.046 0.931 8.5 66.069 ;
    END
  END PAD
  OBS
    LAYER MET1 SPACING 0.09 ;
      RECT 0 -20 65 110 ;
    LAYER MET2 SPACING 0.1 ;
      RECT 62.015 -20 65 110 ;
      RECT 50.83 -20 60.465 110 ;
      RECT 48.245 -20 49.28 110 ;
      RECT 45.685 -20 46.695 110 ;
      RECT 38.41 -20 44.135 110 ;
      RECT 30.245 -20 36.86 110 ;
      RECT 27.315 -20 28.695 110 ;
      RECT 22.77 -20 25.765 110 ;
      RECT 15.56 -20 21.22 110 ;
      RECT 9.7 -20 14.01 110 ;
      RECT 7.025 -20 8.15 110 ;
      RECT 0 -20 5.475 110 ;
      RECT 0 -20 65 109.225 ;
    LAYER MET3 SPACING 0.1 ;
      RECT 0 63.675 65 68.325 ;
      RECT 1.675 -20 65 68.325 ;
      RECT 1.375 63.652 65 68.325 ;
      RECT 1.651 63.387 65 68.325 ;
      RECT 1.421 63.606 65 68.325 ;
      RECT 1.605 63.422 65 68.325 ;
      RECT 1.467 63.56 65 68.325 ;
      RECT 1.559 63.468 65 68.325 ;
      RECT 1.513 63.514 65 68.325 ;
      RECT 1.651 55.887 65 57.613 ;
      RECT 1.605 55.922 65 57.578 ;
      RECT 1.559 55.968 65 57.532 ;
      RECT 1.513 56.014 65 57.486 ;
      RECT 1.467 56.06 65 57.44 ;
      RECT 1.421 56.106 65 57.394 ;
      RECT 1.375 56.152 65 57.348 ;
      RECT 0 56.175 65 57.325 ;
      RECT 1.651 42.387 65 44.113 ;
      RECT 1.605 42.422 65 44.078 ;
      RECT 1.559 42.468 65 44.032 ;
      RECT 1.513 42.514 65 43.986 ;
      RECT 1.467 42.56 65 43.94 ;
      RECT 1.421 42.606 65 43.894 ;
      RECT 1.375 42.652 65 43.848 ;
      RECT 0 42.675 65 43.825 ;
      RECT 1.651 28.887 65 30.613 ;
      RECT 1.605 28.922 65 30.578 ;
      RECT 1.559 28.968 65 30.532 ;
      RECT 1.513 29.014 65 30.486 ;
      RECT 1.467 29.06 65 30.44 ;
      RECT 1.421 29.106 65 30.394 ;
      RECT 1.375 29.152 65 30.348 ;
      RECT 0 29.175 65 30.325 ;
      RECT 1.651 15.387 65 17.113 ;
      RECT 1.605 15.422 65 17.078 ;
      RECT 1.559 15.468 65 17.032 ;
      RECT 1.513 15.514 65 16.986 ;
      RECT 1.467 15.56 65 16.94 ;
      RECT 1.421 15.606 65 16.894 ;
      RECT 1.375 15.652 65 16.848 ;
      RECT 0 15.675 65 16.825 ;
      RECT 1.651 -20 65 3.613 ;
      RECT 1.605 -20 65 3.578 ;
      RECT 1.559 -20 65 3.532 ;
      RECT 1.513 -20 65 3.486 ;
      RECT 1.467 -20 65 3.44 ;
      RECT 1.421 -20 65 3.394 ;
      RECT 1.375 -20 65 3.348 ;
      RECT 0 -20 65 3.325 ;
      RECT 62.015 107.675 65 110 ;
      RECT 50.83 107.675 60.465 110 ;
      RECT 48.245 107.675 49.28 110 ;
      RECT 45.685 107.675 46.695 110 ;
      RECT 38.41 107.675 44.135 110 ;
      RECT 30.245 107.675 36.86 110 ;
      RECT 27.315 107.675 28.695 110 ;
      RECT 22.77 107.675 25.765 110 ;
      RECT 15.56 107.675 21.22 110 ;
      RECT 9.7 107.675 14.01 110 ;
      RECT 7.025 107.675 8.15 110 ;
      RECT 0 107.675 5.475 110 ;
      RECT 0 107.675 65 109.225 ;
      RECT 0 77.175 65 78.325 ;
      RECT 0 89.675 65 90.825 ;
      RECT 0 98.175 65 99.325 ;
    LAYER MET4 SPACING 0.1 ;
      RECT 0 63.675 65 68.325 ;
      RECT 1.675 -20 65 68.325 ;
      RECT 1.375 63.652 65 68.325 ;
      RECT 1.651 63.387 65 68.325 ;
      RECT 1.421 63.606 65 68.325 ;
      RECT 1.605 63.422 65 68.325 ;
      RECT 1.467 63.56 65 68.325 ;
      RECT 1.559 63.468 65 68.325 ;
      RECT 1.513 63.514 65 68.325 ;
      RECT 1.651 55.887 65 57.613 ;
      RECT 1.605 55.922 65 57.578 ;
      RECT 1.559 55.968 65 57.532 ;
      RECT 1.513 56.014 65 57.486 ;
      RECT 1.467 56.06 65 57.44 ;
      RECT 1.421 56.106 65 57.394 ;
      RECT 1.375 56.152 65 57.348 ;
      RECT 0 56.175 65 57.325 ;
      RECT 1.651 42.387 65 44.113 ;
      RECT 1.605 42.422 65 44.078 ;
      RECT 1.559 42.468 65 44.032 ;
      RECT 1.513 42.514 65 43.986 ;
      RECT 1.467 42.56 65 43.94 ;
      RECT 1.421 42.606 65 43.894 ;
      RECT 1.375 42.652 65 43.848 ;
      RECT 0 42.675 65 43.825 ;
      RECT 1.651 28.887 65 30.613 ;
      RECT 1.605 28.922 65 30.578 ;
      RECT 1.559 28.968 65 30.532 ;
      RECT 1.513 29.014 65 30.486 ;
      RECT 1.467 29.06 65 30.44 ;
      RECT 1.421 29.106 65 30.394 ;
      RECT 1.375 29.152 65 30.348 ;
      RECT 0 29.175 65 30.325 ;
      RECT 1.651 15.387 65 17.113 ;
      RECT 1.605 15.422 65 17.078 ;
      RECT 1.559 15.468 65 17.032 ;
      RECT 1.513 15.514 65 16.986 ;
      RECT 1.467 15.56 65 16.94 ;
      RECT 1.421 15.606 65 16.894 ;
      RECT 1.375 15.652 65 16.848 ;
      RECT 0 15.675 65 16.825 ;
      RECT 1.651 -20 65 3.613 ;
      RECT 1.605 -20 65 3.578 ;
      RECT 1.559 -20 65 3.532 ;
      RECT 1.513 -20 65 3.486 ;
      RECT 1.467 -20 65 3.44 ;
      RECT 1.421 -20 65 3.394 ;
      RECT 1.375 -20 65 3.348 ;
      RECT 0 -20 65 3.325 ;
      RECT 62.015 107.675 65 110 ;
      RECT 50.83 107.675 60.465 110 ;
      RECT 48.245 107.675 49.28 110 ;
      RECT 45.685 107.675 46.695 110 ;
      RECT 38.41 107.675 44.135 110 ;
      RECT 30.245 107.675 36.86 110 ;
      RECT 27.315 107.675 28.695 110 ;
      RECT 22.77 107.675 25.765 110 ;
      RECT 15.56 107.675 21.22 110 ;
      RECT 9.7 107.675 14.01 110 ;
      RECT 7.025 107.675 8.15 110 ;
      RECT 0 107.675 5.475 110 ;
      RECT 0 107.675 65 109.225 ;
      RECT 0 77.175 65 78.325 ;
      RECT 0 89.675 65 90.825 ;
      RECT 0 98.175 65 99.325 ;
    LAYER MET5 SPACING 0.1 ;
      RECT 0 63.83 65 68.17 ;
      RECT 1.83 -20 65 68.17 ;
      RECT 1.53 63.807 65 68.17 ;
      RECT 1.806 63.542 65 68.17 ;
      RECT 1.576 63.761 65 68.17 ;
      RECT 1.76 63.577 65 68.17 ;
      RECT 1.622 63.715 65 68.17 ;
      RECT 1.714 63.623 65 68.17 ;
      RECT 1.668 63.669 65 68.17 ;
      RECT 1.806 56.042 65 57.458 ;
      RECT 1.76 56.077 65 57.423 ;
      RECT 1.714 56.123 65 57.377 ;
      RECT 1.668 56.169 65 57.331 ;
      RECT 1.622 56.215 65 57.285 ;
      RECT 1.576 56.261 65 57.239 ;
      RECT 1.53 56.307 65 57.193 ;
      RECT 0 56.33 65 57.17 ;
      RECT 1.806 42.542 65 43.958 ;
      RECT 1.76 42.577 65 43.923 ;
      RECT 1.714 42.623 65 43.877 ;
      RECT 1.668 42.669 65 43.831 ;
      RECT 1.622 42.715 65 43.785 ;
      RECT 1.576 42.761 65 43.739 ;
      RECT 1.53 42.807 65 43.693 ;
      RECT 0 42.83 65 43.67 ;
      RECT 1.806 29.042 65 30.458 ;
      RECT 1.76 29.077 65 30.423 ;
      RECT 1.714 29.123 65 30.377 ;
      RECT 1.668 29.169 65 30.331 ;
      RECT 1.622 29.215 65 30.285 ;
      RECT 1.576 29.261 65 30.239 ;
      RECT 1.53 29.307 65 30.193 ;
      RECT 0 29.33 65 30.17 ;
      RECT 1.806 15.542 65 16.958 ;
      RECT 1.76 15.577 65 16.923 ;
      RECT 1.714 15.623 65 16.877 ;
      RECT 1.668 15.669 65 16.831 ;
      RECT 1.622 15.715 65 16.785 ;
      RECT 1.576 15.761 65 16.739 ;
      RECT 1.53 15.807 65 16.693 ;
      RECT 0 15.83 65 16.67 ;
      RECT 1.806 -20 65 3.458 ;
      RECT 1.76 -20 65 3.423 ;
      RECT 1.714 -20 65 3.377 ;
      RECT 1.668 -20 65 3.331 ;
      RECT 1.622 -20 65 3.285 ;
      RECT 1.576 -20 65 3.239 ;
      RECT 1.53 -20 65 3.193 ;
      RECT 0 -20 65 3.17 ;
      RECT 62.17 107.83 65 110 ;
      RECT 50.985 107.83 60.31 110 ;
      RECT 48.4 107.83 49.125 110 ;
      RECT 45.84 107.83 46.54 110 ;
      RECT 38.565 107.83 43.98 110 ;
      RECT 30.4 107.83 36.705 110 ;
      RECT 27.47 107.83 28.54 110 ;
      RECT 22.925 107.83 25.61 110 ;
      RECT 15.715 107.83 21.065 110 ;
      RECT 9.855 107.83 13.855 110 ;
      RECT 7.18 107.83 7.995 110 ;
      RECT 0 107.83 5.32 110 ;
      RECT 0 107.83 65 109.07 ;
      RECT 0 77.33 65 78.17 ;
      RECT 0 89.83 65 90.67 ;
      RECT 0 98.33 65 99.17 ;
    LAYER T4M2 SPACING 0.4 ;
      RECT 64.584 -20 65 -3.193 ;
      RECT 0 -20 0.428 -3.205 ;
      RECT 64.538 -20 65 -3.239 ;
      RECT 0 -20 0.474 -3.251 ;
      RECT 64.492 -20 65 -3.285 ;
      RECT 0 -20 0.52 -3.297 ;
      RECT 64.446 -20 65 -3.331 ;
      RECT 0 -20 0.566 -3.343 ;
      RECT 64.4 -20 65 -3.377 ;
      RECT 0 -20 0.6 -3.383 ;
      RECT 0 -20 65 -3.4 ;
      RECT 62.44 108.1 65 110 ;
      RECT 51.255 108.1 60.04 110 ;
      RECT 38.835 108.1 43.71 110 ;
      RECT 30.67 108.1 36.435 110 ;
      RECT 27.74 108.1 28.27 110 ;
      RECT 23.195 108.1 25.34 110 ;
      RECT 15.985 108.1 20.795 110 ;
      RECT 10.125 108.1 13.585 110 ;
      RECT 0 108.1 5.05 110 ;
      RECT 0 108.1 65 108.8 ;
    LAYER RDL SPACING 2 ;
      RECT 0 -20 65 -5 ;
      RECT 0 72 65 110 ;
      RECT 3.5 5 61.5 63 ;
  END
END P65_1233_PBMUX

MACRO P65_1233_PWE
  CLASS PAD ;
  ORIGIN 0 20 ;
  FOREIGN P65_1233_PWE 0 -20 ;
  SIZE 130 BY 130 ;
  SYMMETRY X Y R90 ;
  SITE IOSite ;
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA2 ;
    ANTENNAPARTIALCUTAREA 0.0486 LAYER VIA4 ;
    PORT
      LAYER MET5 ;
        RECT 42.755 109.4 43.955 110 ;
      LAYER MET4 ;
        RECT 42.755 109.4 43.955 110 ;
      LAYER MET3 ;
        RECT 42.755 109.4 43.955 110 ;
      LAYER MET2 ;
        RECT 42.755 109.4 43.955 110 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER MET5 ;
        RECT 0 99.5 130 107.5 ;
      LAYER MET4 ;
        RECT 0 99.5 130 107.5 ;
      LAYER MET3 ;
        RECT 0 99.5 130 107.5 ;
      LAYER MET2 ;
        RECT 0 99.5 130 107.5 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET5 ;
        RECT 0 68.5 130 77 ;
        RECT 0 30.788 1.5 42.212 ;
        RECT 0 30.753 1.476 42.247 ;
        RECT 0 30.707 1.43 42.293 ;
        RECT 0 30.661 1.384 42.339 ;
        RECT 0 30.615 1.338 42.385 ;
        RECT 0 30.569 1.292 42.431 ;
        RECT 0 30.523 1.246 42.477 ;
        RECT 0 30.5 1.2 42.5 ;
        RECT 0 44.288 1.5 55.712 ;
        RECT 0 44.253 1.476 55.747 ;
        RECT 0 44.207 1.43 55.793 ;
        RECT 0 44.161 1.384 55.839 ;
        RECT 0 44.115 1.338 55.885 ;
        RECT 0 44.069 1.292 55.931 ;
        RECT 0 44.023 1.246 55.977 ;
        RECT 0 44 1.2 56 ;
        RECT 0 57.788 1.5 63.212 ;
        RECT 0 57.753 1.476 63.247 ;
        RECT 0 57.707 1.43 63.293 ;
        RECT 0 57.661 1.384 63.339 ;
        RECT 0 57.615 1.338 63.385 ;
        RECT 0 57.569 1.292 63.431 ;
        RECT 0 57.523 1.246 63.477 ;
        RECT 0 57.5 1.2 63.5 ;
      LAYER MET4 ;
        RECT 0 68.5 130 77 ;
        RECT 0 30.788 1.5 42.212 ;
        RECT 0 30.753 1.476 42.247 ;
        RECT 0 30.707 1.43 42.293 ;
        RECT 0 30.661 1.384 42.339 ;
        RECT 0 30.615 1.338 42.385 ;
        RECT 0 30.569 1.292 42.431 ;
        RECT 0 30.523 1.246 42.477 ;
        RECT 0 30.5 1.2 42.5 ;
        RECT 0 44.288 1.5 55.712 ;
        RECT 0 44.253 1.476 55.747 ;
        RECT 0 44.207 1.43 55.793 ;
        RECT 0 44.161 1.384 55.839 ;
        RECT 0 44.115 1.338 55.885 ;
        RECT 0 44.069 1.292 55.931 ;
        RECT 0 44.023 1.246 55.977 ;
        RECT 0 44 1.2 56 ;
        RECT 0 57.788 1.5 63.212 ;
        RECT 0 57.753 1.476 63.247 ;
        RECT 0 57.707 1.43 63.293 ;
        RECT 0 57.661 1.384 63.339 ;
        RECT 0 57.615 1.338 63.385 ;
        RECT 0 57.569 1.292 63.431 ;
        RECT 0 57.523 1.246 63.477 ;
        RECT 0 57.5 1.2 63.5 ;
      LAYER MET3 ;
        RECT 0 68.5 130 77 ;
        RECT 0 30.788 1.5 42.212 ;
        RECT 0 30.753 1.476 42.247 ;
        RECT 0 30.707 1.43 42.293 ;
        RECT 0 30.661 1.384 42.339 ;
        RECT 0 30.615 1.338 42.385 ;
        RECT 0 30.569 1.292 42.431 ;
        RECT 0 30.523 1.246 42.477 ;
        RECT 0 30.5 1.2 42.5 ;
        RECT 0 44.288 1.5 55.712 ;
        RECT 0 44.253 1.476 55.747 ;
        RECT 0 44.207 1.43 55.793 ;
        RECT 0 44.161 1.384 55.839 ;
        RECT 0 44.115 1.338 55.885 ;
        RECT 0 44.069 1.292 55.931 ;
        RECT 0 44.023 1.246 55.977 ;
        RECT 0 44 1.2 56 ;
        RECT 0 57.788 1.5 63.212 ;
        RECT 0 57.753 1.476 63.247 ;
        RECT 0 57.707 1.43 63.293 ;
        RECT 0 57.661 1.384 63.339 ;
        RECT 0 57.615 1.338 63.385 ;
        RECT 0 57.569 1.292 63.431 ;
        RECT 0 57.523 1.246 63.477 ;
        RECT 0 57.5 1.2 63.5 ;
      LAYER MET2 ;
        RECT 0 30.5 130 42.5 ;
        RECT 0 57.5 130 63.5 ;
        RECT 0 44 130 56 ;
        RECT 124.615 44 125.815 64.974 ;
        RECT 69.231 57.5 125.807 65.001 ;
        RECT 69.277 57.5 125.761 65.047 ;
        RECT 69.285 57.5 125.715 65.07 ;
        RECT 121.345 44 122.935 65.07 ;
        RECT 116.865 44 118.455 65.07 ;
        RECT 112.385 44 113.975 65.07 ;
        RECT 107.905 44 109.495 65.07 ;
        RECT 103.425 44 105.015 65.07 ;
        RECT 98.945 44 100.535 65.07 ;
        RECT 94.465 44 96.055 65.07 ;
        RECT 89.985 44 91.575 65.07 ;
        RECT 85.505 44 87.095 65.07 ;
        RECT 81.025 44 82.615 65.07 ;
        RECT 76.545 44 78.135 65.07 ;
        RECT 72.065 44 73.655 65.07 ;
        RECT 69.185 44 70.385 64.993 ;
        RECT 69.277 57.5 125.715 65.066 ;
        RECT 69.231 57.5 125.761 65.039 ;
        RECT 59.615 44 60.815 64.974 ;
        RECT 4.231 57.5 60.807 65.001 ;
        RECT 4.277 57.5 60.761 65.047 ;
        RECT 4.285 57.5 60.715 65.07 ;
        RECT 56.345 44 57.935 65.07 ;
        RECT 51.865 44 53.455 65.07 ;
        RECT 47.385 44 48.975 65.07 ;
        RECT 42.905 44 44.495 65.07 ;
        RECT 38.425 44 40.015 65.07 ;
        RECT 33.945 44 35.535 65.07 ;
        RECT 29.465 44 31.055 65.07 ;
        RECT 24.985 44 26.575 65.07 ;
        RECT 20.505 44 22.095 65.07 ;
        RECT 16.025 44 17.615 65.07 ;
        RECT 11.545 44 13.135 65.07 ;
        RECT 7.065 44 8.655 65.07 ;
        RECT 4.185 44 5.385 64.993 ;
        RECT 4.277 57.5 60.715 65.066 ;
        RECT 4.231 57.5 60.761 65.039 ;
        RECT 0 68.5 130 77 ;
    END
  END VDDIO
  PIN VSS
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA2 ;
    ANTENNAPARTIALCUTAREA 12.5388 LAYER VIA4 ;
    PORT
      LAYER MET5 ;
        RECT 0 91 130 98 ;
      LAYER MET4 ;
        RECT 0 91 130 98 ;
      LAYER MET3 ;
        RECT 0 91 130 98 ;
      LAYER MET2 ;
        RECT 0 91 130 98 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA2 ;
    ANTENNAPARTIALCUTAREA 19.5048 LAYER VIA4 ;
    PORT
      LAYER MET5 ;
        RECT 0 78.5 130 89.5 ;
        RECT 0 3.788 1.5 15.212 ;
        RECT 0 3.753 1.476 15.247 ;
        RECT 0 3.707 1.43 15.293 ;
        RECT 0 3.661 1.384 15.339 ;
        RECT 0 3.615 1.338 15.385 ;
        RECT 0 3.569 1.292 15.431 ;
        RECT 0 3.523 1.246 15.477 ;
        RECT 0 3.5 1.2 15.5 ;
        RECT 0 17.288 1.5 28.712 ;
        RECT 0 17.253 1.476 28.747 ;
        RECT 0 17.207 1.43 28.793 ;
        RECT 0 17.161 1.384 28.839 ;
        RECT 0 17.115 1.338 28.885 ;
        RECT 0 17.069 1.292 28.931 ;
        RECT 0 17.023 1.246 28.977 ;
        RECT 0 17 1.2 29 ;
      LAYER MET4 ;
        RECT 0 78.5 130 89.5 ;
        RECT 0 3.788 1.5 15.212 ;
        RECT 0 3.753 1.476 15.247 ;
        RECT 0 3.707 1.43 15.293 ;
        RECT 0 3.661 1.384 15.339 ;
        RECT 0 3.615 1.338 15.385 ;
        RECT 0 3.569 1.292 15.431 ;
        RECT 0 3.523 1.246 15.477 ;
        RECT 0 3.5 1.2 15.5 ;
        RECT 0 17.288 1.5 28.712 ;
        RECT 0 17.253 1.476 28.747 ;
        RECT 0 17.207 1.43 28.793 ;
        RECT 0 17.161 1.384 28.839 ;
        RECT 0 17.115 1.338 28.885 ;
        RECT 0 17.069 1.292 28.931 ;
        RECT 0 17.023 1.246 28.977 ;
        RECT 0 17 1.2 29 ;
      LAYER MET3 ;
        RECT 0 78.5 130 89.5 ;
        RECT 0 3.788 1.5 15.212 ;
        RECT 0 3.753 1.476 15.247 ;
        RECT 0 3.707 1.43 15.293 ;
        RECT 0 3.661 1.384 15.339 ;
        RECT 0 3.615 1.338 15.385 ;
        RECT 0 3.569 1.292 15.431 ;
        RECT 0 3.523 1.246 15.477 ;
        RECT 0 3.5 1.2 15.5 ;
        RECT 0 17.288 1.5 28.712 ;
        RECT 0 17.253 1.476 28.747 ;
        RECT 0 17.207 1.43 28.793 ;
        RECT 0 17.161 1.384 28.839 ;
        RECT 0 17.115 1.338 28.885 ;
        RECT 0 17.069 1.292 28.931 ;
        RECT 0 17.023 1.246 28.977 ;
        RECT 0 17 1.2 29 ;
      LAYER MET2 ;
        RECT 0 17 130 29 ;
        RECT 0 3.5 130 15.5 ;
        RECT 124.805 3.5 125.995 29 ;
        RECT 119.225 3.5 120.415 29 ;
        RECT 113.645 3.5 114.835 29 ;
        RECT 108.065 3.5 109.255 29 ;
        RECT 102.485 3.5 103.675 29 ;
        RECT 96.905 3.5 98.095 29 ;
        RECT 91.325 3.5 92.515 29 ;
        RECT 85.745 3.5 86.935 29 ;
        RECT 80.165 3.5 81.355 29 ;
        RECT 74.585 3.5 75.775 29 ;
        RECT 69.005 3.5 70.195 29 ;
        RECT 59.805 3.5 60.995 29 ;
        RECT 54.225 3.5 55.415 29 ;
        RECT 48.645 3.5 49.835 29 ;
        RECT 43.065 3.5 44.255 29 ;
        RECT 37.485 3.5 38.675 29 ;
        RECT 31.905 3.5 33.095 29 ;
        RECT 26.325 3.5 27.515 29 ;
        RECT 20.745 3.5 21.935 29 ;
        RECT 15.165 3.5 16.355 29 ;
        RECT 9.585 3.5 10.775 29 ;
        RECT 4.005 3.5 5.195 29 ;
        RECT 0 78.5 130 89.5 ;
    END
  END VSSIO
  PIN XC
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA2 ;
    ANTENNAPARTIALCUTAREA 0.0486 LAYER VIA4 ;
    PORT
      LAYER MET5 ;
        RECT 38.275 109.4 39.475 110 ;
      LAYER MET4 ;
        RECT 38.275 109.4 39.475 110 ;
      LAYER MET3 ;
        RECT 38.275 109.4 39.475 110 ;
      LAYER MET2 ;
        RECT 38.275 109.4 39.475 110 ;
    END
  END XC
  PIN XIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER T4M2 ;
        RECT 122 1.08 126.9 66.02 ;
        RECT 122 1.047 126.88 66.053 ;
        RECT 122 1.001 126.834 66.099 ;
        RECT 122 0.955 126.788 66.145 ;
        RECT 122 0.909 126.742 66.191 ;
        RECT 122 0.863 126.696 66.237 ;
        RECT 122 0.817 126.65 66.283 ;
        RECT 122 0.771 126.604 66.329 ;
        RECT 122 0.725 126.558 66.375 ;
        RECT 122 0.679 126.512 66.421 ;
        RECT 122 0.633 126.466 66.467 ;
        RECT 122 0.587 126.42 66.513 ;
        RECT 122 0.541 126.374 66.559 ;
        RECT 122 0.495 126.328 66.605 ;
        RECT 122 0.449 126.282 66.651 ;
        RECT 122 0.403 126.236 66.697 ;
        RECT 122 0.357 126.19 66.743 ;
        RECT 122 0.311 126.144 66.789 ;
        RECT 122 0.265 126.098 66.835 ;
        RECT 122 0.219 126.052 66.881 ;
        RECT 122 0.173 126.006 66.927 ;
        RECT 69.04 57.4 125.96 66.95 ;
        RECT 68.1 43.4 126.9 50.9 ;
        RECT 68.1 29.4 126.9 36.9 ;
        RECT 68.1 15.4 126.9 22.9 ;
        RECT 69.045 0.15 125.96 8.9 ;
        RECT 108 0.15 115.5 66.95 ;
        RECT 94 0.15 101.5 66.95 ;
        RECT 80 0.15 87.5 66.95 ;
        RECT 68.1 1.072 73.5 66.033 ;
        RECT 69.04 0.152 73.5 66.95 ;
        RECT 69.02 0.165 73.5 66.94 ;
        RECT 68.974 0.198 73.5 66.907 ;
        RECT 68.928 0.244 73.5 66.861 ;
        RECT 68.882 0.29 73.5 66.815 ;
        RECT 68.836 0.336 73.5 66.769 ;
        RECT 68.79 0.382 73.5 66.723 ;
        RECT 68.744 0.428 73.5 66.677 ;
        RECT 68.698 0.474 73.5 66.631 ;
        RECT 68.652 0.52 73.5 66.585 ;
        RECT 68.606 0.566 73.5 66.539 ;
        RECT 68.56 0.612 73.5 66.493 ;
        RECT 68.514 0.658 73.5 66.447 ;
        RECT 68.468 0.704 73.5 66.401 ;
        RECT 68.422 0.75 73.5 66.355 ;
        RECT 68.376 0.796 73.5 66.309 ;
        RECT 68.33 0.842 73.5 66.263 ;
        RECT 68.284 0.888 73.5 66.217 ;
        RECT 68.238 0.934 73.5 66.171 ;
        RECT 68.192 0.98 73.5 66.125 ;
        RECT 68.146 1.026 73.5 66.079 ;
    END
  END XIN
  PIN XOUT
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER T4M2 ;
        RECT 57 1.16 61.9 66.02 ;
        RECT 57 1.127 61.88 66.053 ;
        RECT 57 1.081 61.834 66.099 ;
        RECT 57 1.035 61.788 66.145 ;
        RECT 57 0.989 61.742 66.191 ;
        RECT 57 0.943 61.696 66.237 ;
        RECT 57 0.897 61.65 66.283 ;
        RECT 57 0.851 61.604 66.329 ;
        RECT 57 0.805 61.558 66.375 ;
        RECT 57 0.759 61.512 66.421 ;
        RECT 57 0.713 61.466 66.467 ;
        RECT 57 0.667 61.42 66.513 ;
        RECT 57 0.621 61.374 66.559 ;
        RECT 57 0.575 61.328 66.605 ;
        RECT 57 0.529 61.282 66.651 ;
        RECT 57 0.483 61.236 66.697 ;
        RECT 57 0.437 61.19 66.743 ;
        RECT 57 0.391 61.144 66.789 ;
        RECT 57 0.345 61.098 66.835 ;
        RECT 57 0.299 61.052 66.881 ;
        RECT 57 0.253 61.006 66.927 ;
        RECT 4.04 57.355 60.96 66.95 ;
        RECT 57 0.213 60.96 66.95 ;
        RECT 4.132 0.205 60.926 8.855 ;
        RECT 57 0.173 60.926 66.95 ;
        RECT 4.178 0.166 60.88 8.855 ;
        RECT 3.1 43.355 61.9 50.855 ;
        RECT 3.1 29.355 61.9 36.855 ;
        RECT 3.1 15.355 61.9 22.855 ;
        RECT 4.21 0.15 60.88 8.855 ;
        RECT 43 0.15 50.5 66.95 ;
        RECT 29 0.15 36.5 66.95 ;
        RECT 15 0.15 22.5 66.95 ;
        RECT 3.1 1.237 8.5 66.033 ;
        RECT 3.146 1.191 61.9 8.855 ;
        RECT 4.086 0.251 8.5 66.95 ;
        RECT 4.04 0.297 8.5 66.95 ;
        RECT 4.02 0.33 8.5 66.94 ;
        RECT 3.974 0.363 8.5 66.907 ;
        RECT 3.928 0.409 8.5 66.861 ;
        RECT 3.882 0.455 8.5 66.815 ;
        RECT 3.836 0.501 8.5 66.769 ;
        RECT 3.79 0.547 8.5 66.723 ;
        RECT 3.744 0.593 8.5 66.677 ;
        RECT 3.698 0.639 8.5 66.631 ;
        RECT 3.652 0.685 8.5 66.585 ;
        RECT 3.606 0.731 8.5 66.539 ;
        RECT 3.56 0.777 8.5 66.493 ;
        RECT 3.514 0.823 8.5 66.447 ;
        RECT 3.468 0.869 8.5 66.401 ;
        RECT 3.422 0.915 8.5 66.355 ;
        RECT 3.376 0.961 8.5 66.309 ;
        RECT 3.33 1.007 8.5 66.263 ;
        RECT 3.284 1.053 8.5 66.217 ;
        RECT 3.238 1.099 8.5 66.171 ;
        RECT 3.192 1.145 8.5 66.125 ;
        RECT 3.146 57.355 61.834 66.079 ;
    END
  END XOUT
  OBS
    LAYER MET1 SPACING 0.09 ;
      RECT 0 -20 130 110 ;
    LAYER MET2 SPACING 0.1 ;
      RECT 0 65.245 130 68.325 ;
      RECT 125.99 63.675 130 68.325 ;
      RECT 125.89 65.222 130 68.325 ;
      RECT 125.982 65.149 130 68.325 ;
      RECT 60.89 65.241 69.11 68.325 ;
      RECT 0 65.241 4.11 68.325 ;
      RECT 60.89 65.222 69.102 68.325 ;
      RECT 60.936 65.214 69.102 68.325 ;
      RECT 0 65.214 4.102 68.325 ;
      RECT 125.936 65.176 130 68.325 ;
      RECT 60.936 65.176 69.056 68.325 ;
      RECT 60.982 65.168 69.056 68.325 ;
      RECT 0 65.168 4.056 68.325 ;
      RECT 60.982 65.149 69.01 68.325 ;
      RECT 60.99 63.675 69.01 68.325 ;
      RECT 0 63.675 4.01 68.325 ;
      RECT 44.13 107.675 130 110 ;
      RECT 39.65 107.675 42.58 110 ;
      RECT 0 107.675 38.1 110 ;
      RECT 0 107.675 130 109.225 ;
      RECT 0 -20 130 3.325 ;
      RECT 126.17 15.675 130 16.825 ;
      RECT 0 29.175 130 30.325 ;
      RECT 0 42.675 130 43.825 ;
      RECT 125.99 56.175 130 57.325 ;
      RECT 0 77.175 130 78.325 ;
      RECT 0 89.675 130 90.825 ;
      RECT 0 98.175 130 99.325 ;
      RECT 120.59 15.675 124.63 16.825 ;
      RECT 123.11 56.175 124.44 57.325 ;
      RECT 118.63 56.175 121.17 57.325 ;
      RECT 115.01 15.675 119.05 16.825 ;
      RECT 114.15 56.175 116.69 57.325 ;
      RECT 109.43 15.675 113.47 16.825 ;
      RECT 109.67 56.175 112.21 57.325 ;
      RECT 103.85 15.675 107.89 16.825 ;
      RECT 105.19 56.175 107.73 57.325 ;
      RECT 100.71 56.175 103.25 57.325 ;
      RECT 98.27 15.675 102.31 16.825 ;
      RECT 96.23 56.175 98.77 57.325 ;
      RECT 92.69 15.675 96.73 16.825 ;
      RECT 91.75 56.175 94.29 57.325 ;
      RECT 87.11 15.675 91.15 16.825 ;
      RECT 87.27 56.175 89.81 57.325 ;
      RECT 81.53 15.675 85.57 16.825 ;
      RECT 82.79 56.175 85.33 57.325 ;
      RECT 78.31 56.175 80.85 57.325 ;
      RECT 75.95 15.675 79.99 16.825 ;
      RECT 73.83 56.175 76.37 57.325 ;
      RECT 70.37 15.675 74.41 16.825 ;
      RECT 70.56 56.175 71.89 57.325 ;
      RECT 60.99 56.175 69.01 57.325 ;
      RECT 61.17 15.675 68.83 16.825 ;
      RECT 55.59 15.675 59.63 16.825 ;
      RECT 58.11 56.175 59.44 57.325 ;
      RECT 53.63 56.175 56.17 57.325 ;
      RECT 50.01 15.675 54.05 16.825 ;
      RECT 49.15 56.175 51.69 57.325 ;
      RECT 44.43 15.675 48.47 16.825 ;
      RECT 44.67 56.175 47.21 57.325 ;
      RECT 38.85 15.675 42.89 16.825 ;
      RECT 40.19 56.175 42.73 57.325 ;
      RECT 35.71 56.175 38.25 57.325 ;
      RECT 33.27 15.675 37.31 16.825 ;
      RECT 31.23 56.175 33.77 57.325 ;
      RECT 27.69 15.675 31.73 16.825 ;
      RECT 26.75 56.175 29.29 57.325 ;
      RECT 22.11 15.675 26.15 16.825 ;
      RECT 22.27 56.175 24.81 57.325 ;
      RECT 16.53 15.675 20.57 16.825 ;
      RECT 17.79 56.175 20.33 57.325 ;
      RECT 13.31 56.175 15.85 57.325 ;
      RECT 10.95 15.675 14.99 16.825 ;
      RECT 8.83 56.175 11.37 57.325 ;
      RECT 5.37 15.675 9.41 16.825 ;
      RECT 5.56 56.175 6.89 57.325 ;
      RECT 0 56.175 4.01 57.325 ;
      RECT 0 15.675 3.83 16.825 ;
    LAYER MET3 SPACING 0.1 ;
      RECT 0 63.675 130 68.325 ;
      RECT 1.375 63.665 130 68.325 ;
      RECT 68 57.55 127 68.325 ;
      RECT 122 -20 127 68.325 ;
      RECT 3 57.55 62 68.325 ;
      RECT 57 -20 62 68.325 ;
      RECT 108 -20 115.5 68.325 ;
      RECT 94 -20 101.5 68.325 ;
      RECT 80 -20 87.5 68.325 ;
      RECT 68 -20 73.5 68.325 ;
      RECT 43 -20 50.5 68.325 ;
      RECT 29 -20 36.5 68.325 ;
      RECT 15 -20 22.5 68.325 ;
      RECT 3 -20 8.5 68.325 ;
      RECT 122 56.165 130 57.335 ;
      RECT 108 56.165 116.7 57.335 ;
      RECT 91.74 56.165 103.26 57.335 ;
      RECT 78.3 56.165 89.82 57.335 ;
      RECT 57 56.165 73.5 57.335 ;
      RECT 43 56.165 51.7 57.335 ;
      RECT 26.74 56.165 38.26 57.335 ;
      RECT 13.3 56.165 24.82 57.335 ;
      RECT 1.375 56.165 8.5 57.335 ;
      RECT 0 56.175 8.5 57.325 ;
      RECT 68 42.665 127 51.05 ;
      RECT 3 42.665 62 51.05 ;
      RECT 1.375 42.665 130 43.835 ;
      RECT 0 42.675 130 43.825 ;
      RECT 68 29.165 127 37.05 ;
      RECT 3 29.165 62 37.05 ;
      RECT 1.375 29.165 130 30.335 ;
      RECT 0 29.175 130 30.325 ;
      RECT 68 15.55 127 23.05 ;
      RECT 3 15.55 62 23.05 ;
      RECT 1.375 15.665 130 16.835 ;
      RECT 0 15.675 130 16.825 ;
      RECT 68 -20 127 9.05 ;
      RECT 3 -20 62 9.05 ;
      RECT 1.375 -20 130 3.335 ;
      RECT 0 -20 130 3.325 ;
      RECT 128.8 3.5 130 15.5 ;
      RECT 128.776 3.512 130 15.488 ;
      RECT 128.73 3.547 130 15.453 ;
      RECT 128.684 3.593 130 15.407 ;
      RECT 128.638 3.639 130 15.361 ;
      RECT 128.592 3.685 130 15.315 ;
      RECT 128.546 3.731 130 15.269 ;
      RECT 128.5 3.777 130 15.223 ;
      RECT 128.8 17 130 29 ;
      RECT 128.776 17.012 130 28.988 ;
      RECT 128.73 17.047 130 28.953 ;
      RECT 128.684 17.093 130 28.907 ;
      RECT 128.638 17.139 130 28.861 ;
      RECT 128.592 17.185 130 28.815 ;
      RECT 128.546 17.231 130 28.769 ;
      RECT 128.5 17.277 130 28.723 ;
      RECT 128.8 30.5 130 42.5 ;
      RECT 128.776 30.512 130 42.488 ;
      RECT 128.73 30.547 130 42.453 ;
      RECT 128.684 30.593 130 42.407 ;
      RECT 128.638 30.639 130 42.361 ;
      RECT 128.592 30.685 130 42.315 ;
      RECT 128.546 30.731 130 42.269 ;
      RECT 128.5 30.777 130 42.223 ;
      RECT 128.8 44 130 56 ;
      RECT 128.776 44.012 130 55.988 ;
      RECT 128.73 44.047 130 55.953 ;
      RECT 128.684 44.093 130 55.907 ;
      RECT 128.638 44.139 130 55.861 ;
      RECT 128.592 44.185 130 55.815 ;
      RECT 128.546 44.231 130 55.769 ;
      RECT 128.5 44.277 130 55.723 ;
      RECT 128.8 57.5 130 63.5 ;
      RECT 128.776 57.512 130 63.488 ;
      RECT 128.73 57.547 130 63.453 ;
      RECT 128.684 57.593 130 63.407 ;
      RECT 128.638 57.639 130 63.361 ;
      RECT 128.592 57.685 130 63.315 ;
      RECT 128.546 57.731 130 63.269 ;
      RECT 128.5 57.777 130 63.223 ;
      RECT 44.13 107.675 130 110 ;
      RECT 39.65 107.675 42.58 110 ;
      RECT 0 107.675 38.1 110 ;
      RECT 0 107.675 130 109.225 ;
      RECT 63.8 3.5 66.2 15.5 ;
      RECT 63.776 3.512 66.2 15.488 ;
      RECT 63.776 3.523 66.246 15.477 ;
      RECT 63.73 3.547 66.246 15.453 ;
      RECT 63.73 3.569 66.292 15.431 ;
      RECT 63.684 3.593 66.292 15.407 ;
      RECT 63.684 3.615 66.338 15.385 ;
      RECT 63.638 3.639 66.338 15.361 ;
      RECT 63.638 3.661 66.384 15.339 ;
      RECT 63.592 3.685 66.384 15.315 ;
      RECT 63.592 3.707 66.43 15.293 ;
      RECT 63.546 3.731 66.43 15.269 ;
      RECT 63.546 3.753 66.476 15.247 ;
      RECT 63.5 3.777 66.476 15.223 ;
      RECT 63.5 3.788 66.5 15.212 ;
      RECT 63.8 17 66.2 29 ;
      RECT 63.776 17.012 66.2 28.988 ;
      RECT 63.776 17.023 66.246 28.977 ;
      RECT 63.73 17.047 66.246 28.953 ;
      RECT 63.73 17.069 66.292 28.931 ;
      RECT 63.684 17.093 66.292 28.907 ;
      RECT 63.684 17.115 66.338 28.885 ;
      RECT 63.638 17.139 66.338 28.861 ;
      RECT 63.638 17.161 66.384 28.839 ;
      RECT 63.592 17.185 66.384 28.815 ;
      RECT 63.592 17.207 66.43 28.793 ;
      RECT 63.546 17.231 66.43 28.769 ;
      RECT 63.546 17.253 66.476 28.747 ;
      RECT 63.5 17.277 66.476 28.723 ;
      RECT 63.5 17.288 66.5 28.712 ;
      RECT 63.8 30.5 66.2 42.5 ;
      RECT 63.776 30.512 66.2 42.488 ;
      RECT 63.776 30.523 66.246 42.477 ;
      RECT 63.73 30.547 66.246 42.453 ;
      RECT 63.73 30.569 66.292 42.431 ;
      RECT 63.684 30.593 66.292 42.407 ;
      RECT 63.684 30.615 66.338 42.385 ;
      RECT 63.638 30.639 66.338 42.361 ;
      RECT 63.638 30.661 66.384 42.339 ;
      RECT 63.592 30.685 66.384 42.315 ;
      RECT 63.592 30.707 66.43 42.293 ;
      RECT 63.546 30.731 66.43 42.269 ;
      RECT 63.546 30.753 66.476 42.247 ;
      RECT 63.5 30.777 66.476 42.223 ;
      RECT 63.5 30.788 66.5 42.212 ;
      RECT 63.8 44 66.2 56 ;
      RECT 63.776 44.012 66.2 55.988 ;
      RECT 63.776 44.023 66.246 55.977 ;
      RECT 63.73 44.047 66.246 55.953 ;
      RECT 63.73 44.069 66.292 55.931 ;
      RECT 63.684 44.093 66.292 55.907 ;
      RECT 63.684 44.115 66.338 55.885 ;
      RECT 63.638 44.139 66.338 55.861 ;
      RECT 63.638 44.161 66.384 55.839 ;
      RECT 63.592 44.185 66.384 55.815 ;
      RECT 63.592 44.207 66.43 55.793 ;
      RECT 63.546 44.231 66.43 55.769 ;
      RECT 63.546 44.253 66.476 55.747 ;
      RECT 63.5 44.277 66.476 55.723 ;
      RECT 63.5 44.288 66.5 55.712 ;
      RECT 63.8 57.5 66.2 63.5 ;
      RECT 63.776 57.512 66.2 63.488 ;
      RECT 63.776 57.523 66.246 63.477 ;
      RECT 63.73 57.547 66.246 63.453 ;
      RECT 63.73 57.569 66.292 63.431 ;
      RECT 63.684 57.593 66.292 63.407 ;
      RECT 63.684 57.615 66.338 63.385 ;
      RECT 63.638 57.639 66.338 63.361 ;
      RECT 63.638 57.661 66.384 63.339 ;
      RECT 63.592 57.685 66.384 63.315 ;
      RECT 63.592 57.707 66.43 63.293 ;
      RECT 63.546 57.731 66.43 63.269 ;
      RECT 63.546 57.753 66.476 63.247 ;
      RECT 63.5 57.777 66.476 63.223 ;
      RECT 63.5 57.788 66.5 63.212 ;
      RECT 0 77.175 130 78.325 ;
      RECT 0 89.675 130 90.825 ;
      RECT 0 98.175 130 99.325 ;
      RECT 118.62 56.165 121.18 57.335 ;
      RECT 105.18 56.165 107.74 57.335 ;
      RECT 73.82 56.165 76.38 57.335 ;
      RECT 53.62 56.165 56.18 57.335 ;
      RECT 40.18 56.165 42.74 57.335 ;
      RECT 8.82 56.165 11.38 57.335 ;
    LAYER MET4 SPACING 0.1 ;
      RECT 0 63.675 130 68.325 ;
      RECT 1.675 -20 130 68.325 ;
      RECT 1.375 63.652 130 68.325 ;
      RECT 1.651 63.387 130 68.325 ;
      RECT 1.421 63.606 130 68.325 ;
      RECT 1.605 63.422 130 68.325 ;
      RECT 1.467 63.56 130 68.325 ;
      RECT 1.559 63.468 130 68.325 ;
      RECT 1.513 63.514 130 68.325 ;
      RECT 1.651 55.887 130 57.613 ;
      RECT 1.605 55.922 130 57.578 ;
      RECT 1.559 55.968 130 57.532 ;
      RECT 1.513 56.014 130 57.486 ;
      RECT 1.467 56.06 130 57.44 ;
      RECT 1.421 56.106 130 57.394 ;
      RECT 1.375 56.152 130 57.348 ;
      RECT 0 56.175 130 57.325 ;
      RECT 1.651 42.387 130 44.113 ;
      RECT 1.605 42.422 130 44.078 ;
      RECT 1.559 42.468 130 44.032 ;
      RECT 1.513 42.514 130 43.986 ;
      RECT 1.467 42.56 130 43.94 ;
      RECT 1.421 42.606 130 43.894 ;
      RECT 1.375 42.652 130 43.848 ;
      RECT 0 42.675 130 43.825 ;
      RECT 1.651 28.887 130 30.613 ;
      RECT 1.605 28.922 130 30.578 ;
      RECT 1.559 28.968 130 30.532 ;
      RECT 1.513 29.014 130 30.486 ;
      RECT 1.467 29.06 130 30.44 ;
      RECT 1.421 29.106 130 30.394 ;
      RECT 1.375 29.152 130 30.348 ;
      RECT 0 29.175 130 30.325 ;
      RECT 1.651 15.387 130 17.113 ;
      RECT 1.605 15.422 130 17.078 ;
      RECT 1.559 15.468 130 17.032 ;
      RECT 1.513 15.514 130 16.986 ;
      RECT 1.467 15.56 130 16.94 ;
      RECT 1.421 15.606 130 16.894 ;
      RECT 1.375 15.652 130 16.848 ;
      RECT 0 15.675 130 16.825 ;
      RECT 1.651 -20 130 3.613 ;
      RECT 1.605 -20 130 3.578 ;
      RECT 1.559 -20 130 3.532 ;
      RECT 1.513 -20 130 3.486 ;
      RECT 1.467 -20 130 3.44 ;
      RECT 1.421 -20 130 3.394 ;
      RECT 1.375 -20 130 3.348 ;
      RECT 0 -20 130 3.325 ;
      RECT 44.13 107.675 130 110 ;
      RECT 39.65 107.675 42.58 110 ;
      RECT 0 107.675 38.1 110 ;
      RECT 0 107.675 130 109.225 ;
      RECT 0 77.175 130 78.325 ;
      RECT 0 89.675 130 90.825 ;
      RECT 0 98.175 130 99.325 ;
    LAYER MET5 SPACING 0.1 ;
      RECT 0 63.83 130 68.17 ;
      RECT 1.83 -20 130 68.17 ;
      RECT 1.53 63.807 130 68.17 ;
      RECT 1.806 63.542 130 68.17 ;
      RECT 1.576 63.761 130 68.17 ;
      RECT 1.76 63.577 130 68.17 ;
      RECT 1.622 63.715 130 68.17 ;
      RECT 1.714 63.623 130 68.17 ;
      RECT 1.668 63.669 130 68.17 ;
      RECT 1.806 56.042 130 57.458 ;
      RECT 1.76 56.077 130 57.423 ;
      RECT 1.714 56.123 130 57.377 ;
      RECT 1.668 56.169 130 57.331 ;
      RECT 1.622 56.215 130 57.285 ;
      RECT 1.576 56.261 130 57.239 ;
      RECT 1.53 56.307 130 57.193 ;
      RECT 0 56.33 130 57.17 ;
      RECT 1.806 42.542 130 43.958 ;
      RECT 1.76 42.577 130 43.923 ;
      RECT 1.714 42.623 130 43.877 ;
      RECT 1.668 42.669 130 43.831 ;
      RECT 1.622 42.715 130 43.785 ;
      RECT 1.576 42.761 130 43.739 ;
      RECT 1.53 42.807 130 43.693 ;
      RECT 0 42.83 130 43.67 ;
      RECT 1.806 29.042 130 30.458 ;
      RECT 1.76 29.077 130 30.423 ;
      RECT 1.714 29.123 130 30.377 ;
      RECT 1.668 29.169 130 30.331 ;
      RECT 1.622 29.215 130 30.285 ;
      RECT 1.576 29.261 130 30.239 ;
      RECT 1.53 29.307 130 30.193 ;
      RECT 0 29.33 130 30.17 ;
      RECT 1.806 15.542 130 16.958 ;
      RECT 1.76 15.577 130 16.923 ;
      RECT 1.714 15.623 130 16.877 ;
      RECT 1.668 15.669 130 16.831 ;
      RECT 1.622 15.715 130 16.785 ;
      RECT 1.576 15.761 130 16.739 ;
      RECT 1.53 15.807 130 16.693 ;
      RECT 0 15.83 130 16.67 ;
      RECT 1.806 -20 130 3.458 ;
      RECT 1.76 -20 130 3.423 ;
      RECT 1.714 -20 130 3.377 ;
      RECT 1.668 -20 130 3.331 ;
      RECT 1.622 -20 130 3.285 ;
      RECT 1.576 -20 130 3.239 ;
      RECT 1.53 -20 130 3.193 ;
      RECT 0 -20 130 3.17 ;
      RECT 44.285 107.83 130 110 ;
      RECT 39.805 107.83 42.425 110 ;
      RECT 0 107.83 37.945 110 ;
      RECT 0 107.83 130 109.07 ;
      RECT 0 77.33 130 78.17 ;
      RECT 0 89.83 130 90.67 ;
      RECT 0 98.33 130 99.17 ;
    LAYER T4M2 SPACING 0.4 ;
      RECT 64.728 -20 65.16 -2.779 ;
      RECT 64.728 -20 65.206 -2.788 ;
      RECT 64.682 -20 65.206 -2.825 ;
      RECT 64.682 -20 65.252 -2.834 ;
      RECT 0 -20 0.436 -2.853 ;
      RECT 64.636 -20 65.252 -2.871 ;
      RECT 64.636 -20 65.298 -2.88 ;
      RECT 0 -20 0.482 -2.899 ;
      RECT 64.59 -20 65.298 -2.917 ;
      RECT 64.59 -20 65.344 -2.926 ;
      RECT 0 -20 0.528 -2.945 ;
      RECT 64.544 -20 65.344 -2.963 ;
      RECT 64.544 -20 65.39 -2.972 ;
      RECT 0 -20 0.574 -2.991 ;
      RECT 129.59 -20 130 -2.997 ;
      RECT 64.498 -20 65.39 -3.009 ;
      RECT 64.498 -20 65.436 -3.018 ;
      RECT 0 -20 0.62 -3.037 ;
      RECT 129.544 -20 130 -3.043 ;
      RECT 64.452 -20 65.436 -3.055 ;
      RECT 64.452 -20 65.482 -3.064 ;
      RECT 0 -20 0.64 -3.07 ;
      RECT 129.498 -20 130 -3.089 ;
      RECT 64.406 -20 65.482 -3.101 ;
      RECT 0 -20 0.686 -3.103 ;
      RECT 64.406 -20 65.528 -3.11 ;
      RECT 129.452 -20 130 -3.135 ;
      RECT 64.36 -20 65.528 -3.147 ;
      RECT 0 -20 0.732 -3.149 ;
      RECT 64.36 -20 65.574 -3.156 ;
      RECT 129.406 -20 130 -3.181 ;
      RECT 64.326 -20 65.574 -3.187 ;
      RECT 0 -20 0.778 -3.195 ;
      RECT 64.326 -20 65.62 -3.202 ;
      RECT 129.36 -20 130 -3.227 ;
      RECT 64.28 -20 65.62 -3.227 ;
      RECT 0 -20 0.81 -3.234 ;
      RECT 64.28 -20 65.64 -3.235 ;
      RECT 64.28 -20 65.645 -3.248 ;
      RECT 0 -20 130 -3.25 ;
      RECT 44.555 108.1 130 110 ;
      RECT 40.075 108.1 42.155 110 ;
      RECT 0 108.1 37.675 110 ;
      RECT 0 108.1 130 108.8 ;
    LAYER RDL SPACING 2 ;
      RECT 0 -20 130 -4.85 ;
      RECT 0 71.95 130 110 ;
      RECT 68 4.5 127 63.5 ;
      RECT 3 4.5 62 63.5 ;
  END
END P65_1233_PWE

MACRO P65_1233_VDD1
  CLASS PAD ;
  ORIGIN 0 20 ;
  FOREIGN P65_1233_VDD1 0 -20 ;
  SIZE 65 BY 130 ;
  SYMMETRY X Y R90 ;
  SITE IOSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET2 ;
        RECT 0 99.98 6.5 107.02 ;
        RECT 0 99.937 6.46 107.063 ;
        RECT 0 99.891 6.414 107.109 ;
        RECT 0 99.845 6.368 107.155 ;
        RECT 0 99.799 6.322 107.201 ;
        RECT 0 99.753 6.276 107.247 ;
        RECT 0 99.707 6.23 107.293 ;
        RECT 0 99.661 6.184 107.339 ;
        RECT 0 99.615 6.138 107.385 ;
        RECT 0 99.569 6.092 107.431 ;
        RECT 0 99.523 6.046 107.477 ;
        RECT 0 99.5 6 107.5 ;
    END
    PORT
      CLASS CORE ;
      LAYER MET5 ;
        RECT 0 99.5 65 107.5 ;
      LAYER MET4 ;
        RECT 0 99.5 65 107.5 ;
      LAYER MET3 ;
        RECT 0 99.5 65 107.5 ;
    END
  END VDD
  PIN VDD1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET5 ;
        RECT 8 109 57 110 ;
      LAYER T4M2 ;
        RECT 57 4.532 61.9 65.968 ;
        RECT 57 4.497 61.875 66.003 ;
        RECT 57 4.451 61.829 66.049 ;
        RECT 57 4.405 61.783 66.095 ;
        RECT 57 4.359 61.737 66.141 ;
        RECT 57 4.313 61.691 66.187 ;
        RECT 57 4.267 61.645 66.233 ;
        RECT 57 4.221 61.599 66.279 ;
        RECT 57 4.175 61.553 66.325 ;
        RECT 57 4.129 61.507 66.371 ;
        RECT 57 4.083 61.461 66.417 ;
        RECT 57 4.037 61.415 66.463 ;
        RECT 57 3.991 61.369 66.509 ;
        RECT 57 3.945 61.323 66.555 ;
        RECT 57 3.899 61.277 66.601 ;
        RECT 57 3.853 61.231 66.647 ;
        RECT 57 3.807 61.185 66.693 ;
        RECT 57 3.761 61.139 66.739 ;
        RECT 57 3.715 61.093 66.785 ;
        RECT 57 3.669 61.047 66.831 ;
        RECT 57 3.623 61.001 66.877 ;
        RECT 4.045 57.5 60.955 66.9 ;
        RECT 57 3.595 60.955 66.9 ;
        RECT 4.045 3.577 60.946 9 ;
        RECT 57 3.568 60.946 66.9 ;
        RECT 4.091 3.549 60.9 9 ;
        RECT 3.1 43.5 61.9 51 ;
        RECT 3.1 29.5 61.9 37 ;
        RECT 3.1 15.5 61.9 23 ;
        RECT 4.1 0.1 60.9 9 ;
        RECT 43 0.1 50.5 66.9 ;
        RECT 29 0.1 36.5 66.9 ;
        RECT 15 0.1 22.5 66.9 ;
        RECT 3.1 4.522 8.5 65.978 ;
        RECT 4.02 3.612 8.5 66.888 ;
        RECT 3.974 3.648 8.5 66.852 ;
        RECT 3.928 3.694 8.5 66.806 ;
        RECT 3.882 3.74 8.5 66.76 ;
        RECT 3.836 3.786 8.5 66.714 ;
        RECT 3.79 3.832 8.5 66.668 ;
        RECT 3.744 3.878 8.5 66.622 ;
        RECT 3.698 3.924 8.5 66.576 ;
        RECT 3.652 3.97 8.5 66.53 ;
        RECT 3.606 4.016 8.5 66.484 ;
        RECT 3.56 4.062 8.5 66.438 ;
        RECT 3.514 4.108 8.5 66.392 ;
        RECT 3.468 4.154 8.5 66.346 ;
        RECT 3.422 4.2 8.5 66.3 ;
        RECT 3.376 4.246 8.5 66.254 ;
        RECT 3.33 4.292 8.5 66.208 ;
        RECT 3.284 4.338 8.5 66.162 ;
        RECT 3.238 4.384 8.5 66.116 ;
        RECT 3.192 4.43 8.5 66.07 ;
        RECT 3.146 4.476 8.5 66.024 ;
      LAYER MET4 ;
        RECT 8 109 57 110 ;
      LAYER MET3 ;
        RECT 8 109 57 110 ;
      LAYER MET2 ;
        RECT 8 99.5 57 110 ;
        RECT 45.92 78.5 57 110 ;
        RECT 8 78.5 57 89.5 ;
        RECT 33.32 78.5 44.32 110 ;
        RECT 20.66 78.5 31.66 110 ;
        RECT 8 78.5 19 110 ;
    END
  END VDD1
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET5 ;
        RECT 0 68.5 65 77 ;
        RECT 0 30.788 1.5 42.212 ;
        RECT 0 30.753 1.476 42.247 ;
        RECT 0 30.707 1.43 42.293 ;
        RECT 0 30.661 1.384 42.339 ;
        RECT 0 30.615 1.338 42.385 ;
        RECT 0 30.569 1.292 42.431 ;
        RECT 0 30.523 1.246 42.477 ;
        RECT 0 30.5 1.2 42.5 ;
        RECT 0 44.288 1.5 55.712 ;
        RECT 0 44.253 1.476 55.747 ;
        RECT 0 44.207 1.43 55.793 ;
        RECT 0 44.161 1.384 55.839 ;
        RECT 0 44.115 1.338 55.885 ;
        RECT 0 44.069 1.292 55.931 ;
        RECT 0 44.023 1.246 55.977 ;
        RECT 0 44 1.2 56 ;
        RECT 0 57.788 1.5 63.212 ;
        RECT 0 57.753 1.476 63.247 ;
        RECT 0 57.707 1.43 63.293 ;
        RECT 0 57.661 1.384 63.339 ;
        RECT 0 57.615 1.338 63.385 ;
        RECT 0 57.569 1.292 63.431 ;
        RECT 0 57.523 1.246 63.477 ;
        RECT 0 57.5 1.2 63.5 ;
      LAYER MET4 ;
        RECT 0 68.5 65 77 ;
        RECT 0 30.788 1.5 42.212 ;
        RECT 0 30.753 1.476 42.247 ;
        RECT 0 30.707 1.43 42.293 ;
        RECT 0 30.661 1.384 42.339 ;
        RECT 0 30.615 1.338 42.385 ;
        RECT 0 30.569 1.292 42.431 ;
        RECT 0 30.523 1.246 42.477 ;
        RECT 0 30.5 1.2 42.5 ;
        RECT 0 44.288 1.5 55.712 ;
        RECT 0 44.253 1.476 55.747 ;
        RECT 0 44.207 1.43 55.793 ;
        RECT 0 44.161 1.384 55.839 ;
        RECT 0 44.115 1.338 55.885 ;
        RECT 0 44.069 1.292 55.931 ;
        RECT 0 44.023 1.246 55.977 ;
        RECT 0 44 1.2 56 ;
        RECT 0 57.788 1.5 63.212 ;
        RECT 0 57.753 1.476 63.247 ;
        RECT 0 57.707 1.43 63.293 ;
        RECT 0 57.661 1.384 63.339 ;
        RECT 0 57.615 1.338 63.385 ;
        RECT 0 57.569 1.292 63.431 ;
        RECT 0 57.523 1.246 63.477 ;
        RECT 0 57.5 1.2 63.5 ;
      LAYER MET3 ;
        RECT 0 68.5 65 77 ;
        RECT 0 30.788 1.5 42.212 ;
        RECT 0 30.753 1.476 42.247 ;
        RECT 0 30.707 1.43 42.293 ;
        RECT 0 30.661 1.384 42.339 ;
        RECT 0 30.615 1.338 42.385 ;
        RECT 0 30.569 1.292 42.431 ;
        RECT 0 30.523 1.246 42.477 ;
        RECT 0 30.5 1.2 42.5 ;
        RECT 0 44.288 1.5 55.712 ;
        RECT 0 44.253 1.476 55.747 ;
        RECT 0 44.207 1.43 55.793 ;
        RECT 0 44.161 1.384 55.839 ;
        RECT 0 44.115 1.338 55.885 ;
        RECT 0 44.069 1.292 55.931 ;
        RECT 0 44.023 1.246 55.977 ;
        RECT 0 44 1.2 56 ;
        RECT 0 57.788 1.5 63.212 ;
        RECT 0 57.753 1.476 63.247 ;
        RECT 0 57.707 1.43 63.293 ;
        RECT 0 57.661 1.384 63.339 ;
        RECT 0 57.615 1.338 63.385 ;
        RECT 0 57.569 1.292 63.431 ;
        RECT 0 57.523 1.246 63.477 ;
        RECT 0 57.5 1.2 63.5 ;
      LAYER MET2 ;
        RECT 0 68.5 65 77 ;
        RECT 0 57.5 65 63.5 ;
        RECT 0 44 65 56 ;
        RECT 0 30.5 65 42.5 ;
        RECT 57.015 30.5 58.205 77 ;
        RECT 51.435 30.5 52.625 77 ;
        RECT 45.855 30.5 47.045 77 ;
        RECT 40.275 30.5 41.465 77 ;
        RECT 34.695 30.5 35.885 77 ;
        RECT 29.115 30.5 30.305 77 ;
        RECT 23.535 30.5 24.725 77 ;
        RECT 17.955 30.5 19.145 77 ;
        RECT 12.375 30.5 13.565 77 ;
        RECT 6.795 30.5 7.985 77 ;
    END
  END VDDIO
  PIN VSS
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 6.2694 LAYER VIA4 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 1.6848 LAYER VIA2 ;
    PORT
      LAYER MET5 ;
        RECT 0 91 65 98 ;
      LAYER MET4 ;
        RECT 0 91 65 98 ;
      LAYER MET3 ;
        RECT 0 91 65 98 ;
      LAYER MET2 ;
        RECT 0 91.48 6.5 97.52 ;
        RECT 0 91.437 6.46 97.563 ;
        RECT 0 91.391 6.414 97.609 ;
        RECT 0 91.345 6.368 97.655 ;
        RECT 0 91.299 6.322 97.701 ;
        RECT 0 91.253 6.276 97.747 ;
        RECT 0 91.207 6.23 97.793 ;
        RECT 0 91.161 6.184 97.839 ;
        RECT 0 91.115 6.138 97.885 ;
        RECT 0 91.069 6.092 97.931 ;
        RECT 0 91.023 6.046 97.977 ;
        RECT 0 91 6 98 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA2 ;
    ANTENNAPARTIALCUTAREA 9.7524 LAYER VIA4 ;
    PORT
      LAYER MET5 ;
        RECT 0 78.5 65 89.5 ;
        RECT 0 3.788 1.5 15.212 ;
        RECT 0 3.753 1.476 15.247 ;
        RECT 0 3.707 1.43 15.293 ;
        RECT 0 3.661 1.384 15.339 ;
        RECT 0 3.615 1.338 15.385 ;
        RECT 0 3.569 1.292 15.431 ;
        RECT 0 3.523 1.246 15.477 ;
        RECT 0 3.5 1.2 15.5 ;
        RECT 0 17.288 1.5 28.712 ;
        RECT 0 17.253 1.476 28.747 ;
        RECT 0 17.207 1.43 28.793 ;
        RECT 0 17.161 1.384 28.839 ;
        RECT 0 17.115 1.338 28.885 ;
        RECT 0 17.069 1.292 28.931 ;
        RECT 0 17.023 1.246 28.977 ;
        RECT 0 17 1.2 29 ;
      LAYER MET4 ;
        RECT 0 78.5 65 89.5 ;
        RECT 0 3.788 1.5 15.212 ;
        RECT 0 3.753 1.476 15.247 ;
        RECT 0 3.707 1.43 15.293 ;
        RECT 0 3.661 1.384 15.339 ;
        RECT 0 3.615 1.338 15.385 ;
        RECT 0 3.569 1.292 15.431 ;
        RECT 0 3.523 1.246 15.477 ;
        RECT 0 3.5 1.2 15.5 ;
        RECT 0 17.288 1.5 28.712 ;
        RECT 0 17.253 1.476 28.747 ;
        RECT 0 17.207 1.43 28.793 ;
        RECT 0 17.161 1.384 28.839 ;
        RECT 0 17.115 1.338 28.885 ;
        RECT 0 17.069 1.292 28.931 ;
        RECT 0 17.023 1.246 28.977 ;
        RECT 0 17 1.2 29 ;
      LAYER MET3 ;
        RECT 0 78.5 65 89.5 ;
        RECT 0 3.788 1.5 15.212 ;
        RECT 0 3.753 1.476 15.247 ;
        RECT 0 3.707 1.43 15.293 ;
        RECT 0 3.661 1.384 15.339 ;
        RECT 0 3.615 1.338 15.385 ;
        RECT 0 3.569 1.292 15.431 ;
        RECT 0 3.523 1.246 15.477 ;
        RECT 0 3.5 1.2 15.5 ;
        RECT 0 17.288 1.5 28.712 ;
        RECT 0 17.253 1.476 28.747 ;
        RECT 0 17.207 1.43 28.793 ;
        RECT 0 17.161 1.384 28.839 ;
        RECT 0 17.115 1.338 28.885 ;
        RECT 0 17.069 1.292 28.931 ;
        RECT 0 17.023 1.246 28.977 ;
        RECT 0 17 1.2 29 ;
      LAYER MET2 ;
        RECT 0 17 65 29 ;
        RECT 0 3.5 65 15.5 ;
        RECT 59.805 3.5 60.995 29 ;
        RECT 54.225 3.5 55.415 29 ;
        RECT 48.645 3.5 49.835 29 ;
        RECT 43.065 3.5 44.255 29 ;
        RECT 37.485 3.5 38.675 29 ;
        RECT 31.905 3.5 33.095 29 ;
        RECT 26.325 3.5 27.515 29 ;
        RECT 20.745 3.5 21.935 29 ;
        RECT 15.165 3.5 16.355 29 ;
        RECT 9.585 3.5 10.775 29 ;
        RECT 4.005 3.5 5.195 29 ;
        RECT 0 78.98 6.5 89.02 ;
        RECT 0 78.937 6.46 89.063 ;
        RECT 0 78.891 6.414 89.109 ;
        RECT 0 78.845 6.368 89.155 ;
        RECT 0 78.799 6.322 89.201 ;
        RECT 0 78.753 6.276 89.247 ;
        RECT 0 78.707 6.23 89.293 ;
        RECT 0 78.661 6.184 89.339 ;
        RECT 0 78.615 6.138 89.385 ;
        RECT 0 78.569 6.092 89.431 ;
        RECT 0 78.523 6.046 89.477 ;
        RECT 0 78.5 6 89.5 ;
    END
  END VSSIO
  OBS
    LAYER MET1 SPACING 0.09 ;
      RECT 0 -20 65 110 ;
    LAYER MET2 SPACING 0.1 ;
      RECT 57.175 77.175 65 110 ;
      RECT 0 107.675 7.825 110 ;
      RECT 6.675 77.175 7.825 110 ;
      RECT 6.175 107.652 7.825 110 ;
      RECT 6.635 107.195 7.825 110 ;
      RECT 6.221 107.606 7.825 110 ;
      RECT 6.589 107.238 7.825 110 ;
      RECT 6.267 107.56 7.825 110 ;
      RECT 6.543 107.284 7.825 110 ;
      RECT 6.313 107.514 7.825 110 ;
      RECT 6.497 107.33 7.825 110 ;
      RECT 6.359 107.468 7.825 110 ;
      RECT 6.451 107.376 7.825 110 ;
      RECT 6.405 107.422 7.825 110 ;
      RECT 6.635 97.695 7.825 99.805 ;
      RECT 6.589 97.738 7.825 99.762 ;
      RECT 6.543 97.784 7.825 99.716 ;
      RECT 6.497 97.83 7.825 99.67 ;
      RECT 6.451 97.876 7.825 99.624 ;
      RECT 6.405 97.922 7.825 99.578 ;
      RECT 6.359 97.968 7.825 99.532 ;
      RECT 6.313 98.014 7.825 99.486 ;
      RECT 6.267 98.06 7.825 99.44 ;
      RECT 6.221 98.106 7.825 99.394 ;
      RECT 6.175 98.152 7.825 99.348 ;
      RECT 0 98.175 7.825 99.325 ;
      RECT 6.635 89.195 7.825 91.305 ;
      RECT 6.589 89.238 7.825 91.262 ;
      RECT 6.543 89.284 7.825 91.216 ;
      RECT 6.497 89.33 7.825 91.17 ;
      RECT 6.451 89.376 7.825 91.124 ;
      RECT 6.405 89.422 7.825 91.078 ;
      RECT 6.359 89.468 7.825 91.032 ;
      RECT 6.313 89.514 7.825 90.986 ;
      RECT 6.267 89.56 7.825 90.94 ;
      RECT 6.221 89.606 7.825 90.894 ;
      RECT 6.175 89.652 7.825 90.848 ;
      RECT 0 89.675 7.825 90.825 ;
      RECT 6.635 77.175 7.825 78.805 ;
      RECT 6.589 77.175 7.825 78.762 ;
      RECT 6.543 77.175 7.825 78.716 ;
      RECT 6.497 77.175 7.825 78.67 ;
      RECT 6.451 77.175 7.825 78.624 ;
      RECT 6.405 77.175 7.825 78.578 ;
      RECT 6.359 77.175 7.825 78.532 ;
      RECT 6.313 77.175 7.825 78.486 ;
      RECT 6.267 77.175 7.825 78.44 ;
      RECT 6.221 77.175 7.825 78.394 ;
      RECT 6.175 77.175 7.825 78.348 ;
      RECT 0 77.175 65 78.325 ;
      RECT 0 -20 65 3.325 ;
      RECT 61.17 15.675 65 16.825 ;
      RECT 0 29.175 65 30.325 ;
      RECT 58.38 42.675 65 43.825 ;
      RECT 58.38 56.175 65 57.325 ;
      RECT 58.38 63.675 65 68.325 ;
      RECT 55.59 15.675 59.63 16.825 ;
      RECT 52.8 42.675 56.84 43.825 ;
      RECT 52.8 56.175 56.84 57.325 ;
      RECT 52.8 63.675 56.84 68.325 ;
      RECT 50.01 15.675 54.05 16.825 ;
      RECT 47.22 42.675 51.26 43.825 ;
      RECT 47.22 56.175 51.26 57.325 ;
      RECT 47.22 63.675 51.26 68.325 ;
      RECT 44.43 15.675 48.47 16.825 ;
      RECT 44.495 89.675 45.745 99.325 ;
      RECT 41.64 42.675 45.68 43.825 ;
      RECT 41.64 56.175 45.68 57.325 ;
      RECT 41.64 63.675 45.68 68.325 ;
      RECT 38.85 15.675 42.89 16.825 ;
      RECT 36.06 42.675 40.1 43.825 ;
      RECT 36.06 56.175 40.1 57.325 ;
      RECT 36.06 63.675 40.1 68.325 ;
      RECT 33.27 15.675 37.31 16.825 ;
      RECT 30.48 42.675 34.52 43.825 ;
      RECT 30.48 56.175 34.52 57.325 ;
      RECT 30.48 63.675 34.52 68.325 ;
      RECT 31.835 89.675 33.145 99.325 ;
      RECT 27.69 15.675 31.73 16.825 ;
      RECT 24.9 42.675 28.94 43.825 ;
      RECT 24.9 56.175 28.94 57.325 ;
      RECT 24.9 63.675 28.94 68.325 ;
      RECT 22.11 15.675 26.15 16.825 ;
      RECT 19.32 42.675 23.36 43.825 ;
      RECT 19.32 56.175 23.36 57.325 ;
      RECT 19.32 63.675 23.36 68.325 ;
      RECT 16.53 15.675 20.57 16.825 ;
      RECT 19.175 89.675 20.485 99.325 ;
      RECT 13.74 42.675 17.78 43.825 ;
      RECT 13.74 56.175 17.78 57.325 ;
      RECT 13.74 63.675 17.78 68.325 ;
      RECT 10.95 15.675 14.99 16.825 ;
      RECT 8.16 42.675 12.2 43.825 ;
      RECT 8.16 56.175 12.2 57.325 ;
      RECT 8.16 63.675 12.2 68.325 ;
      RECT 5.37 15.675 9.41 16.825 ;
      RECT 0 42.675 6.62 43.825 ;
      RECT 0 56.175 6.62 57.325 ;
      RECT 0 63.675 6.62 68.325 ;
      RECT 0 15.675 3.83 16.825 ;
    LAYER MET3 SPACING 0.1 ;
      RECT 62 63.665 65 68.325 ;
      RECT 58.37 -20 61 68.325 ;
      RECT 52.79 57.5 56.85 68.325 ;
      RECT 47.21 57.5 51.27 68.325 ;
      RECT 41.63 57.5 45.69 68.325 ;
      RECT 36.05 57.5 40.11 68.325 ;
      RECT 30.47 -20 34.53 68.325 ;
      RECT 24.89 57.5 28.95 68.325 ;
      RECT 19.31 57.5 23.37 68.325 ;
      RECT 13.73 57.5 17.79 68.325 ;
      RECT 8.15 57.5 12.21 68.325 ;
      RECT 4 -20 6.63 68.325 ;
      RECT 0 63.675 3 68.325 ;
      RECT 1.375 63.665 3 68.325 ;
      RECT 4 57.5 61 67 ;
      RECT 57 -20 61 67 ;
      RECT 43 -20 50.5 67 ;
      RECT 29 -20 36.5 67 ;
      RECT 15 -20 22.5 67 ;
      RECT 4 -20 8.5 67 ;
      RECT 62 56.165 65 57.335 ;
      RECT 41.63 56.165 51.27 57.335 ;
      RECT 24.89 56.165 40.11 57.335 ;
      RECT 13.73 56.165 23.37 57.335 ;
      RECT 4 56.165 12.21 57.335 ;
      RECT 1.375 56.165 3 57.335 ;
      RECT 0 56.175 3 57.325 ;
      RECT 4 43.5 61 51 ;
      RECT 62 42.665 65 43.835 ;
      RECT 1.375 42.665 3 43.835 ;
      RECT 0 42.675 3 43.825 ;
      RECT 52.79 42.665 56.85 51 ;
      RECT 41.63 42.665 51.27 51 ;
      RECT 24.89 42.665 40.11 51 ;
      RECT 13.73 42.665 23.37 51 ;
      RECT 4 42.665 12.21 51 ;
      RECT 4 29.165 61 37 ;
      RECT 62 29.165 65 30.335 ;
      RECT 1.375 29.165 3 30.335 ;
      RECT 0 29.175 3 30.325 ;
      RECT 4 15.5 61 23 ;
      RECT 62 15.665 65 16.835 ;
      RECT 1.375 15.665 3 16.835 ;
      RECT 0 15.675 3 16.825 ;
      RECT 4 -20 61 9 ;
      RECT 1.375 -20 65 3.335 ;
      RECT 0 -20 65 3.325 ;
      RECT 61.966 4.483 62 68.325 ;
      RECT 61.92 4.443 61.966 68.325 ;
      RECT 61.874 4.397 61.92 68.325 ;
      RECT 61.828 4.351 61.874 68.325 ;
      RECT 61.782 4.305 61.828 68.325 ;
      RECT 61.736 4.259 61.782 68.325 ;
      RECT 61.69 4.213 61.736 68.325 ;
      RECT 61.644 4.167 61.69 68.325 ;
      RECT 61.598 4.121 61.644 68.325 ;
      RECT 61.552 4.075 61.598 68.325 ;
      RECT 61.506 4.029 61.552 68.325 ;
      RECT 61.46 3.983 61.506 68.325 ;
      RECT 61.414 3.937 61.46 68.325 ;
      RECT 61.368 3.891 61.414 68.325 ;
      RECT 61.322 3.845 61.368 68.325 ;
      RECT 61.276 3.799 61.322 68.325 ;
      RECT 61.23 3.753 61.276 68.325 ;
      RECT 61.184 3.707 61.23 68.325 ;
      RECT 61.138 3.661 61.184 68.325 ;
      RECT 61.092 3.615 61.138 68.325 ;
      RECT 61.046 3.569 61.092 68.325 ;
      RECT 61 3.523 61.046 68.325 ;
      RECT 3.966 3.517 4 68.325 ;
      RECT 3.92 3.557 3.966 68.325 ;
      RECT 3.874 3.603 3.92 68.325 ;
      RECT 3.828 3.649 3.874 68.325 ;
      RECT 3.782 3.695 3.828 68.325 ;
      RECT 3.736 3.741 3.782 68.325 ;
      RECT 3.69 3.787 3.736 68.325 ;
      RECT 3.644 3.833 3.69 68.325 ;
      RECT 3.598 3.879 3.644 68.325 ;
      RECT 3.552 3.925 3.598 68.325 ;
      RECT 3.506 3.971 3.552 68.325 ;
      RECT 3.46 4.017 3.506 68.325 ;
      RECT 3.414 4.063 3.46 68.325 ;
      RECT 3.368 4.109 3.414 68.325 ;
      RECT 3.322 4.155 3.368 68.325 ;
      RECT 3.276 4.201 3.322 68.325 ;
      RECT 3.23 4.247 3.276 68.325 ;
      RECT 3.184 4.293 3.23 68.325 ;
      RECT 3.138 4.339 3.184 68.325 ;
      RECT 3.092 4.385 3.138 68.325 ;
      RECT 3.046 4.431 3.092 68.325 ;
      RECT 3 4.477 3.046 68.325 ;
      RECT 63.8 3.5 65 15.5 ;
      RECT 63.776 3.512 65 15.488 ;
      RECT 63.73 3.547 65 15.453 ;
      RECT 63.684 3.593 65 15.407 ;
      RECT 63.638 3.639 65 15.361 ;
      RECT 63.592 3.685 65 15.315 ;
      RECT 63.546 3.731 65 15.269 ;
      RECT 63.5 3.777 65 15.223 ;
      RECT 63.8 17 65 29 ;
      RECT 63.776 17.012 65 28.988 ;
      RECT 63.73 17.047 65 28.953 ;
      RECT 63.684 17.093 65 28.907 ;
      RECT 63.638 17.139 65 28.861 ;
      RECT 63.592 17.185 65 28.815 ;
      RECT 63.546 17.231 65 28.769 ;
      RECT 63.5 17.277 65 28.723 ;
      RECT 63.8 30.5 65 42.5 ;
      RECT 63.776 30.512 65 42.488 ;
      RECT 63.73 30.547 65 42.453 ;
      RECT 63.684 30.593 65 42.407 ;
      RECT 63.638 30.639 65 42.361 ;
      RECT 63.592 30.685 65 42.315 ;
      RECT 63.546 30.731 65 42.269 ;
      RECT 63.5 30.777 65 42.223 ;
      RECT 63.8 44 65 56 ;
      RECT 63.776 44.012 65 55.988 ;
      RECT 63.73 44.047 65 55.953 ;
      RECT 63.684 44.093 65 55.907 ;
      RECT 63.638 44.139 65 55.861 ;
      RECT 63.592 44.185 65 55.815 ;
      RECT 63.546 44.231 65 55.769 ;
      RECT 63.5 44.277 65 55.723 ;
      RECT 63.8 57.5 65 63.5 ;
      RECT 63.776 57.512 65 63.488 ;
      RECT 63.73 57.547 65 63.453 ;
      RECT 63.684 57.593 65 63.407 ;
      RECT 63.638 57.639 65 63.361 ;
      RECT 63.592 57.685 65 63.315 ;
      RECT 63.546 57.731 65 63.269 ;
      RECT 63.5 57.777 65 63.223 ;
      RECT 57.175 107.675 65 110 ;
      RECT 57.165 107.675 65 108.825 ;
      RECT 0 107.675 7.825 110 ;
      RECT 0 107.675 7.835 108.825 ;
      RECT 0 77.175 65 78.325 ;
      RECT 57.165 89.675 65 90.825 ;
      RECT 57.165 98.175 65 99.325 ;
      RECT 52.79 56.165 56.85 57.335 ;
      RECT 44.485 89.675 45.755 90.825 ;
      RECT 44.485 98.175 45.755 99.325 ;
      RECT 31.825 89.675 33.155 90.825 ;
      RECT 31.825 98.175 33.155 99.325 ;
      RECT 19.165 89.675 20.495 90.825 ;
      RECT 19.165 98.175 20.495 99.325 ;
      RECT 0 89.675 7.835 90.825 ;
      RECT 0 98.175 7.835 99.325 ;
    LAYER MET4 SPACING 0.1 ;
      RECT 0 63.675 65 68.325 ;
      RECT 1.675 -20 65 68.325 ;
      RECT 1.375 63.652 65 68.325 ;
      RECT 1.651 63.387 65 68.325 ;
      RECT 1.421 63.606 65 68.325 ;
      RECT 1.605 63.422 65 68.325 ;
      RECT 1.467 63.56 65 68.325 ;
      RECT 1.559 63.468 65 68.325 ;
      RECT 1.513 63.514 65 68.325 ;
      RECT 1.651 55.887 65 57.613 ;
      RECT 1.605 55.922 65 57.578 ;
      RECT 1.559 55.968 65 57.532 ;
      RECT 1.513 56.014 65 57.486 ;
      RECT 1.467 56.06 65 57.44 ;
      RECT 1.421 56.106 65 57.394 ;
      RECT 1.375 56.152 65 57.348 ;
      RECT 0 56.175 65 57.325 ;
      RECT 1.651 42.387 65 44.113 ;
      RECT 1.605 42.422 65 44.078 ;
      RECT 1.559 42.468 65 44.032 ;
      RECT 1.513 42.514 65 43.986 ;
      RECT 1.467 42.56 65 43.94 ;
      RECT 1.421 42.606 65 43.894 ;
      RECT 1.375 42.652 65 43.848 ;
      RECT 0 42.675 65 43.825 ;
      RECT 1.651 28.887 65 30.613 ;
      RECT 1.605 28.922 65 30.578 ;
      RECT 1.559 28.968 65 30.532 ;
      RECT 1.513 29.014 65 30.486 ;
      RECT 1.467 29.06 65 30.44 ;
      RECT 1.421 29.106 65 30.394 ;
      RECT 1.375 29.152 65 30.348 ;
      RECT 0 29.175 65 30.325 ;
      RECT 1.651 15.387 65 17.113 ;
      RECT 1.605 15.422 65 17.078 ;
      RECT 1.559 15.468 65 17.032 ;
      RECT 1.513 15.514 65 16.986 ;
      RECT 1.467 15.56 65 16.94 ;
      RECT 1.421 15.606 65 16.894 ;
      RECT 1.375 15.652 65 16.848 ;
      RECT 0 15.675 65 16.825 ;
      RECT 1.651 -20 65 3.613 ;
      RECT 1.605 -20 65 3.578 ;
      RECT 1.559 -20 65 3.532 ;
      RECT 1.513 -20 65 3.486 ;
      RECT 1.467 -20 65 3.44 ;
      RECT 1.421 -20 65 3.394 ;
      RECT 1.375 -20 65 3.348 ;
      RECT 0 -20 65 3.325 ;
      RECT 57.175 107.675 65 110 ;
      RECT 0 107.675 7.825 110 ;
      RECT 0 107.675 65 108.825 ;
      RECT 0 77.175 65 78.325 ;
      RECT 0 89.675 65 90.825 ;
      RECT 0 98.175 65 99.325 ;
    LAYER MET5 SPACING 0.1 ;
      RECT 0 63.83 65 68.17 ;
      RECT 1.83 -20 65 68.17 ;
      RECT 1.53 63.807 65 68.17 ;
      RECT 1.806 63.542 65 68.17 ;
      RECT 1.576 63.761 65 68.17 ;
      RECT 1.76 63.577 65 68.17 ;
      RECT 1.622 63.715 65 68.17 ;
      RECT 1.714 63.623 65 68.17 ;
      RECT 1.668 63.669 65 68.17 ;
      RECT 1.806 56.042 65 57.458 ;
      RECT 1.76 56.077 65 57.423 ;
      RECT 1.714 56.123 65 57.377 ;
      RECT 1.668 56.169 65 57.331 ;
      RECT 1.622 56.215 65 57.285 ;
      RECT 1.576 56.261 65 57.239 ;
      RECT 1.53 56.307 65 57.193 ;
      RECT 0 56.33 65 57.17 ;
      RECT 1.806 42.542 65 43.958 ;
      RECT 1.76 42.577 65 43.923 ;
      RECT 1.714 42.623 65 43.877 ;
      RECT 1.668 42.669 65 43.831 ;
      RECT 1.622 42.715 65 43.785 ;
      RECT 1.576 42.761 65 43.739 ;
      RECT 1.53 42.807 65 43.693 ;
      RECT 0 42.83 65 43.67 ;
      RECT 1.806 29.042 65 30.458 ;
      RECT 1.76 29.077 65 30.423 ;
      RECT 1.714 29.123 65 30.377 ;
      RECT 1.668 29.169 65 30.331 ;
      RECT 1.622 29.215 65 30.285 ;
      RECT 1.576 29.261 65 30.239 ;
      RECT 1.53 29.307 65 30.193 ;
      RECT 0 29.33 65 30.17 ;
      RECT 1.806 15.542 65 16.958 ;
      RECT 1.76 15.577 65 16.923 ;
      RECT 1.714 15.623 65 16.877 ;
      RECT 1.668 15.669 65 16.831 ;
      RECT 1.622 15.715 65 16.785 ;
      RECT 1.576 15.761 65 16.739 ;
      RECT 1.53 15.807 65 16.693 ;
      RECT 0 15.83 65 16.67 ;
      RECT 1.806 -20 65 3.458 ;
      RECT 1.76 -20 65 3.423 ;
      RECT 1.714 -20 65 3.377 ;
      RECT 1.668 -20 65 3.331 ;
      RECT 1.622 -20 65 3.285 ;
      RECT 1.576 -20 65 3.239 ;
      RECT 1.53 -20 65 3.193 ;
      RECT 0 -20 65 3.17 ;
      RECT 57.33 107.83 65 110 ;
      RECT 0 107.83 7.67 110 ;
      RECT 0 107.83 65 108.67 ;
      RECT 0 77.33 65 78.17 ;
      RECT 0 89.83 65 90.67 ;
      RECT 0 98.33 65 99.17 ;
    LAYER T4M2 SPACING 0.4 ;
      RECT 64.585 -20 65 0.453 ;
      RECT 0 -20 0.436 0.432 ;
      RECT 64.539 -20 65 0.407 ;
      RECT 0 -20 0.482 0.386 ;
      RECT 64.493 -20 65 0.361 ;
      RECT 0 -20 0.528 0.34 ;
      RECT 64.447 -20 65 0.315 ;
      RECT 0 -20 0.574 0.294 ;
      RECT 64.401 -20 65 0.269 ;
      RECT 0 -20 0.62 0.248 ;
      RECT 64.355 -20 65 0.223 ;
      RECT 0 -20 0.645 0.212 ;
      RECT 64.346 -20 65 0.195 ;
      RECT 0 -20 0.691 0.177 ;
      RECT 64.3 -20 65 0.168 ;
      RECT 0 -20 0.7 0.149 ;
      RECT 0 -20 65 -3.3 ;
      RECT 57.6 108.1 65 110 ;
      RECT 0 108.1 7.4 110 ;
    LAYER RDL SPACING 2 ;
      RECT 0 -20 65 -4.9 ;
      RECT 0 71.9 65 110 ;
      RECT 3 4.5 62 63.5 ;
  END
END P65_1233_VDD1

MACRO P65_1233_VDD1A
  CLASS PAD ;
  ORIGIN 0 20 ;
  FOREIGN P65_1233_VDD1A 0 -20 ;
  SIZE 65 BY 130 ;
  SYMMETRY X Y R90 ;
  SITE IOSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET4 ;
        RECT 0 100.483 6.5 106.517 ;
        RECT 0 100.443 6.466 106.557 ;
        RECT 0 100.397 6.42 106.603 ;
        RECT 0 100.351 6.374 106.649 ;
        RECT 0 100.305 6.328 106.695 ;
        RECT 0 100.259 6.282 106.741 ;
        RECT 0 100.213 6.236 106.787 ;
        RECT 0 100.167 6.19 106.833 ;
        RECT 0 100.121 6.144 106.879 ;
        RECT 0 100.075 6.098 106.925 ;
        RECT 0 100.029 6.052 106.971 ;
        RECT 0 99.983 6.006 107.017 ;
        RECT 0 99.937 5.96 107.063 ;
        RECT 0 99.891 5.914 107.109 ;
        RECT 0 99.845 5.868 107.155 ;
        RECT 0 99.799 5.822 107.201 ;
        RECT 0 99.753 5.776 107.247 ;
        RECT 0 99.707 5.73 107.293 ;
        RECT 0 99.661 5.684 107.339 ;
        RECT 0 99.615 5.638 107.385 ;
        RECT 0 99.569 5.592 107.431 ;
        RECT 0 99.523 5.546 107.477 ;
        RECT 0 99.5 5.5 107.5 ;
      LAYER MET3 ;
        RECT 0 100.483 6.5 106.517 ;
        RECT 0 100.443 6.466 106.557 ;
        RECT 0 100.397 6.42 106.603 ;
        RECT 0 100.351 6.374 106.649 ;
        RECT 0 100.305 6.328 106.695 ;
        RECT 0 100.259 6.282 106.741 ;
        RECT 0 100.213 6.236 106.787 ;
        RECT 0 100.167 6.19 106.833 ;
        RECT 0 100.121 6.144 106.879 ;
        RECT 0 100.075 6.098 106.925 ;
        RECT 0 100.029 6.052 106.971 ;
        RECT 0 99.983 6.006 107.017 ;
        RECT 0 99.937 5.96 107.063 ;
        RECT 0 99.891 5.914 107.109 ;
        RECT 0 99.845 5.868 107.155 ;
        RECT 0 99.799 5.822 107.201 ;
        RECT 0 99.753 5.776 107.247 ;
        RECT 0 99.707 5.73 107.293 ;
        RECT 0 99.661 5.684 107.339 ;
        RECT 0 99.615 5.638 107.385 ;
        RECT 0 99.569 5.592 107.431 ;
        RECT 0 99.523 5.546 107.477 ;
        RECT 0 99.5 5.5 107.5 ;
    END
    PORT
      CLASS CORE ;
      LAYER MET5 ;
        RECT 0 99.5 65 107.5 ;
      LAYER MET2 ;
        RECT 0 99.5 65 107.5 ;
    END
  END VDD
  PIN VDDA1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET5 ;
        RECT 8 109 57 110 ;
      LAYER T4M2 ;
        RECT 3 68.5 62 77 ;
        RECT 57 4.483 62 63.5 ;
        RECT 57 4.443 61.966 63.5 ;
        RECT 3.046 4.431 61.92 9 ;
        RECT 57 4.397 61.92 63.5 ;
        RECT 3.092 4.385 61.874 9 ;
        RECT 57 4.351 61.874 63.5 ;
        RECT 3.138 4.339 61.828 9 ;
        RECT 57 4.305 61.828 63.5 ;
        RECT 3.184 4.293 61.782 9 ;
        RECT 57 4.259 61.782 63.5 ;
        RECT 3.23 4.247 61.736 9 ;
        RECT 57 4.213 61.736 63.5 ;
        RECT 3.276 4.201 61.69 9 ;
        RECT 57 4.167 61.69 63.5 ;
        RECT 3.322 4.155 61.644 9 ;
        RECT 57 4.121 61.644 63.5 ;
        RECT 3.368 4.109 61.598 9 ;
        RECT 57 4.075 61.598 63.5 ;
        RECT 3.414 4.063 61.552 9 ;
        RECT 57 4.029 61.552 63.5 ;
        RECT 3.46 4.017 61.506 9 ;
        RECT 57 3.983 61.506 63.5 ;
        RECT 3.506 3.971 61.46 9 ;
        RECT 57 3.937 61.46 63.5 ;
        RECT 3.552 3.925 61.414 9 ;
        RECT 57 3.891 61.414 63.5 ;
        RECT 3.598 3.879 61.368 9 ;
        RECT 57 3.845 61.368 63.5 ;
        RECT 3.644 3.833 61.322 9 ;
        RECT 57 3.799 61.322 63.5 ;
        RECT 3.69 3.787 61.276 9 ;
        RECT 57 3.753 61.276 63.5 ;
        RECT 3.736 3.741 61.23 9 ;
        RECT 57 3.707 61.23 63.5 ;
        RECT 3.782 3.695 61.184 9 ;
        RECT 57 3.661 61.184 63.5 ;
        RECT 3.828 3.649 61.138 9 ;
        RECT 57 3.615 61.138 63.5 ;
        RECT 3.874 3.603 61.092 9 ;
        RECT 57 3.569 61.092 63.5 ;
        RECT 3.92 3.557 61.046 9 ;
        RECT 57 3.523 61.046 63.5 ;
        RECT 3.966 3.517 61 9 ;
        RECT 46 57.5 57 77 ;
        RECT 3 43.5 62 51 ;
        RECT 3 29.5 62 37 ;
        RECT 3 15.5 62 23 ;
        RECT 4 0 61 9 ;
        RECT 43 0 50.5 63.5 ;
        RECT 33.27 57.5 44.34 77 ;
        RECT 29 0 36.5 63.5 ;
        RECT 20.66 57.5 31.66 77 ;
        RECT 15 0 22.5 63.5 ;
        RECT 8 57.5 19 77 ;
        RECT 3 4.477 8.5 63.5 ;
      LAYER MET4 ;
        RECT 3 68.5 62 77 ;
        RECT 57 4.483 62 63.5 ;
        RECT 57 4.443 61.966 63.5 ;
        RECT 3.046 4.431 61.92 9 ;
        RECT 57 4.397 61.92 63.5 ;
        RECT 3.092 4.385 61.874 9 ;
        RECT 57 4.351 61.874 63.5 ;
        RECT 3.138 4.339 61.828 9 ;
        RECT 57 4.305 61.828 63.5 ;
        RECT 3.184 4.293 61.782 9 ;
        RECT 57 4.259 61.782 63.5 ;
        RECT 3.23 4.247 61.736 9 ;
        RECT 57 4.213 61.736 63.5 ;
        RECT 3.276 4.201 61.69 9 ;
        RECT 57 4.167 61.69 63.5 ;
        RECT 3.322 4.155 61.644 9 ;
        RECT 57 4.121 61.644 63.5 ;
        RECT 3.368 4.109 61.598 9 ;
        RECT 57 4.075 61.598 63.5 ;
        RECT 3.414 4.063 61.552 9 ;
        RECT 57 4.029 61.552 63.5 ;
        RECT 3.46 4.017 61.506 9 ;
        RECT 57 3.983 61.506 63.5 ;
        RECT 3.506 3.971 61.46 9 ;
        RECT 57 3.937 61.46 63.5 ;
        RECT 3.552 3.925 61.414 9 ;
        RECT 57 3.891 61.414 63.5 ;
        RECT 3.598 3.879 61.368 9 ;
        RECT 57 3.845 61.368 63.5 ;
        RECT 3.644 3.833 61.322 9 ;
        RECT 57 3.799 61.322 63.5 ;
        RECT 3.69 3.787 61.276 9 ;
        RECT 57 3.753 61.276 63.5 ;
        RECT 3.736 3.741 61.23 9 ;
        RECT 57 3.707 61.23 63.5 ;
        RECT 3.782 3.695 61.184 9 ;
        RECT 57 3.661 61.184 63.5 ;
        RECT 3.828 3.649 61.138 9 ;
        RECT 57 3.615 61.138 63.5 ;
        RECT 3.874 3.603 61.092 9 ;
        RECT 57 3.569 61.092 63.5 ;
        RECT 3.92 3.557 61.046 9 ;
        RECT 57 3.523 61.046 63.5 ;
        RECT 3.966 3.517 61 9 ;
        RECT 8 109 57 110 ;
        RECT 46 57.5 57 110 ;
        RECT 3 43.5 62 51 ;
        RECT 3 29.5 62 37 ;
        RECT 3 15.5 62 23 ;
        RECT 4 0 61 9 ;
        RECT 43 0 50.5 63.5 ;
        RECT 33.27 57.5 44.34 110 ;
        RECT 29 0 36.5 63.5 ;
        RECT 20.66 57.5 31.66 110 ;
        RECT 15 0 22.5 63.5 ;
        RECT 8 57.5 19 110 ;
        RECT 3 4.477 8.5 63.5 ;
      LAYER MET3 ;
        RECT 3 68.5 62 77 ;
        RECT 57 4.483 62 63.5 ;
        RECT 57 4.443 61.966 63.5 ;
        RECT 3.046 4.431 61.92 9 ;
        RECT 57 4.397 61.92 63.5 ;
        RECT 3.092 4.385 61.874 9 ;
        RECT 57 4.351 61.874 63.5 ;
        RECT 3.138 4.339 61.828 9 ;
        RECT 57 4.305 61.828 63.5 ;
        RECT 3.184 4.293 61.782 9 ;
        RECT 57 4.259 61.782 63.5 ;
        RECT 3.23 4.247 61.736 9 ;
        RECT 57 4.213 61.736 63.5 ;
        RECT 3.276 4.201 61.69 9 ;
        RECT 57 4.167 61.69 63.5 ;
        RECT 3.322 4.155 61.644 9 ;
        RECT 57 4.121 61.644 63.5 ;
        RECT 3.368 4.109 61.598 9 ;
        RECT 57 4.075 61.598 63.5 ;
        RECT 3.414 4.063 61.552 9 ;
        RECT 57 4.029 61.552 63.5 ;
        RECT 3.46 4.017 61.506 9 ;
        RECT 57 3.983 61.506 63.5 ;
        RECT 3.506 3.971 61.46 9 ;
        RECT 57 3.937 61.46 63.5 ;
        RECT 3.552 3.925 61.414 9 ;
        RECT 57 3.891 61.414 63.5 ;
        RECT 3.598 3.879 61.368 9 ;
        RECT 57 3.845 61.368 63.5 ;
        RECT 3.644 3.833 61.322 9 ;
        RECT 57 3.799 61.322 63.5 ;
        RECT 3.69 3.787 61.276 9 ;
        RECT 57 3.753 61.276 63.5 ;
        RECT 3.736 3.741 61.23 9 ;
        RECT 57 3.707 61.23 63.5 ;
        RECT 3.782 3.695 61.184 9 ;
        RECT 57 3.661 61.184 63.5 ;
        RECT 3.828 3.649 61.138 9 ;
        RECT 57 3.615 61.138 63.5 ;
        RECT 3.874 3.603 61.092 9 ;
        RECT 57 3.569 61.092 63.5 ;
        RECT 3.92 3.557 61.046 9 ;
        RECT 57 3.523 61.046 63.5 ;
        RECT 3.966 3.517 61 9 ;
        RECT 8 109 57 110 ;
        RECT 46 57.5 57 110 ;
        RECT 3 43.5 62 51 ;
        RECT 3 29.5 62 37 ;
        RECT 3 15.5 62 23 ;
        RECT 4 0 61 9 ;
        RECT 43 0 50.5 63.5 ;
        RECT 33.27 57.5 44.34 110 ;
        RECT 29 0 36.5 63.5 ;
        RECT 20.66 57.5 31.66 110 ;
        RECT 15 0 22.5 63.5 ;
        RECT 8 57.5 19 110 ;
        RECT 3 4.477 8.5 63.5 ;
      LAYER MET2 ;
        RECT 8 109 57 110 ;
    END
  END VDDA1
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET5 ;
        RECT 0 30.788 1.5 42.212 ;
        RECT 0 30.753 1.476 42.247 ;
        RECT 0 30.707 1.43 42.293 ;
        RECT 0 30.661 1.384 42.339 ;
        RECT 0 30.615 1.338 42.385 ;
        RECT 0 30.569 1.292 42.431 ;
        RECT 0 30.523 1.246 42.477 ;
        RECT 0 30.5 1.2 42.5 ;
        RECT 0 44.288 1.5 55.712 ;
        RECT 0 44.253 1.476 55.747 ;
        RECT 0 44.207 1.43 55.793 ;
        RECT 0 44.161 1.384 55.839 ;
        RECT 0 44.115 1.338 55.885 ;
        RECT 0 44.069 1.292 55.931 ;
        RECT 0 44.023 1.246 55.977 ;
        RECT 0 44 1.2 56 ;
        RECT 0 57.788 1.5 63.212 ;
        RECT 0 57.753 1.476 63.247 ;
        RECT 0 57.707 1.43 63.293 ;
        RECT 0 57.661 1.384 63.339 ;
        RECT 0 57.615 1.338 63.385 ;
        RECT 0 57.569 1.292 63.431 ;
        RECT 0 57.523 1.246 63.477 ;
        RECT 0 57.5 1.2 63.5 ;
        RECT 0 68.788 1.5 76.712 ;
        RECT 0 68.753 1.476 76.747 ;
        RECT 0 68.707 1.43 76.793 ;
        RECT 0 68.661 1.384 76.839 ;
        RECT 0 68.615 1.338 76.885 ;
        RECT 0 68.569 1.292 76.931 ;
        RECT 0 68.523 1.246 76.977 ;
        RECT 0 68.5 1.2 77 ;
      LAYER MET4 ;
        RECT 0 30.788 1.5 42.212 ;
        RECT 0 30.753 1.476 42.247 ;
        RECT 0 30.707 1.43 42.293 ;
        RECT 0 30.661 1.384 42.339 ;
        RECT 0 30.615 1.338 42.385 ;
        RECT 0 30.569 1.292 42.431 ;
        RECT 0 30.523 1.246 42.477 ;
        RECT 0 30.5 1.2 42.5 ;
        RECT 0 44.288 1.5 55.712 ;
        RECT 0 44.253 1.476 55.747 ;
        RECT 0 44.207 1.43 55.793 ;
        RECT 0 44.161 1.384 55.839 ;
        RECT 0 44.115 1.338 55.885 ;
        RECT 0 44.069 1.292 55.931 ;
        RECT 0 44.023 1.246 55.977 ;
        RECT 0 44 1.2 56 ;
        RECT 0 57.788 1.5 63.212 ;
        RECT 0 57.753 1.476 63.247 ;
        RECT 0 57.707 1.43 63.293 ;
        RECT 0 57.661 1.384 63.339 ;
        RECT 0 57.615 1.338 63.385 ;
        RECT 0 57.569 1.292 63.431 ;
        RECT 0 57.523 1.246 63.477 ;
        RECT 0 57.5 1.2 63.5 ;
        RECT 0 68.788 1.5 76.712 ;
        RECT 0 68.753 1.476 76.747 ;
        RECT 0 68.707 1.43 76.793 ;
        RECT 0 68.661 1.384 76.839 ;
        RECT 0 68.615 1.338 76.885 ;
        RECT 0 68.569 1.292 76.931 ;
        RECT 0 68.523 1.246 76.977 ;
        RECT 0 68.5 1.2 77 ;
      LAYER MET3 ;
        RECT 0 30.788 1.5 42.212 ;
        RECT 0 30.753 1.476 42.247 ;
        RECT 0 30.707 1.43 42.293 ;
        RECT 0 30.661 1.384 42.339 ;
        RECT 0 30.615 1.338 42.385 ;
        RECT 0 30.569 1.292 42.431 ;
        RECT 0 30.523 1.246 42.477 ;
        RECT 0 30.5 1.2 42.5 ;
        RECT 0 44.288 1.5 55.712 ;
        RECT 0 44.253 1.476 55.747 ;
        RECT 0 44.207 1.43 55.793 ;
        RECT 0 44.161 1.384 55.839 ;
        RECT 0 44.115 1.338 55.885 ;
        RECT 0 44.069 1.292 55.931 ;
        RECT 0 44.023 1.246 55.977 ;
        RECT 0 44 1.2 56 ;
        RECT 0 57.788 1.5 63.212 ;
        RECT 0 57.753 1.476 63.247 ;
        RECT 0 57.707 1.43 63.293 ;
        RECT 0 57.661 1.384 63.339 ;
        RECT 0 57.615 1.338 63.385 ;
        RECT 0 57.569 1.292 63.431 ;
        RECT 0 57.523 1.246 63.477 ;
        RECT 0 57.5 1.2 63.5 ;
        RECT 0 68.788 1.5 76.712 ;
        RECT 0 68.753 1.476 76.747 ;
        RECT 0 68.707 1.43 76.793 ;
        RECT 0 68.661 1.384 76.839 ;
        RECT 0 68.615 1.338 76.885 ;
        RECT 0 68.569 1.292 76.931 ;
        RECT 0 68.523 1.246 76.977 ;
        RECT 0 68.5 1.2 77 ;
      LAYER MET2 ;
        RECT 0 57.5 65 63.5 ;
        RECT 0 44 65 56 ;
        RECT 0 30.5 65 42.5 ;
        RECT 56.015 30.5 59.205 63.5 ;
        RECT 50.435 30.5 53.625 63.5 ;
        RECT 44.855 30.5 48.045 63.5 ;
        RECT 39.275 30.5 42.465 63.5 ;
        RECT 33.695 30.5 36.885 63.5 ;
        RECT 28.115 30.5 31.305 63.5 ;
        RECT 22.535 30.5 25.725 63.5 ;
        RECT 16.955 30.5 20.145 63.5 ;
        RECT 11.375 30.5 14.565 63.5 ;
        RECT 5.795 30.5 8.985 63.5 ;
        RECT 0 68.5 65 77 ;
    END
  END VDDA
  PIN VSS
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 44.5 LAYER MET4 ;
    ANTENNAPARTIALMETALAREA 44.5 LAYER MET3 ;
    ANTENNAPARTIALCUTAREA 1.0692 LAYER VIA4 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 4.617 LAYER VIA2 ;
    PORT
      LAYER MET5 ;
        RECT 0 91 65 98 ;
      LAYER MET4 ;
        RECT 0 91.983 6.5 97.017 ;
        RECT 0 91.943 6.466 97.057 ;
        RECT 0 91.897 6.42 97.103 ;
        RECT 0 91.851 6.374 97.149 ;
        RECT 0 91.805 6.328 97.195 ;
        RECT 0 91.759 6.282 97.241 ;
        RECT 0 91.713 6.236 97.287 ;
        RECT 0 91.667 6.19 97.333 ;
        RECT 0 91.621 6.144 97.379 ;
        RECT 0 91.575 6.098 97.425 ;
        RECT 0 91.529 6.052 97.471 ;
        RECT 0 91.483 6.006 97.517 ;
        RECT 0 91.437 5.96 97.563 ;
        RECT 0 91.391 5.914 97.609 ;
        RECT 0 91.345 5.868 97.655 ;
        RECT 0 91.299 5.822 97.701 ;
        RECT 0 91.253 5.776 97.747 ;
        RECT 0 91.207 5.73 97.793 ;
        RECT 0 91.161 5.684 97.839 ;
        RECT 0 91.115 5.638 97.885 ;
        RECT 0 91.069 5.592 97.931 ;
        RECT 0 91.023 5.546 97.977 ;
        RECT 0 91 5.5 98 ;
      LAYER MET3 ;
        RECT 0 91.983 6.5 97.017 ;
        RECT 0 91.943 6.466 97.057 ;
        RECT 0 91.897 6.42 97.103 ;
        RECT 0 91.851 6.374 97.149 ;
        RECT 0 91.805 6.328 97.195 ;
        RECT 0 91.759 6.282 97.241 ;
        RECT 0 91.713 6.236 97.287 ;
        RECT 0 91.667 6.19 97.333 ;
        RECT 0 91.621 6.144 97.379 ;
        RECT 0 91.575 6.098 97.425 ;
        RECT 0 91.529 6.052 97.471 ;
        RECT 0 91.483 6.006 97.517 ;
        RECT 0 91.437 5.96 97.563 ;
        RECT 0 91.391 5.914 97.609 ;
        RECT 0 91.345 5.868 97.655 ;
        RECT 0 91.299 5.822 97.701 ;
        RECT 0 91.253 5.776 97.747 ;
        RECT 0 91.207 5.73 97.793 ;
        RECT 0 91.161 5.684 97.839 ;
        RECT 0 91.115 5.638 97.885 ;
        RECT 0 91.069 5.592 97.931 ;
        RECT 0 91.023 5.546 97.977 ;
        RECT 0 91 5.5 98 ;
      LAYER MET2 ;
        RECT 0 91 65 98 ;
    END
  END VSS
  PIN VSSA
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 70.5 LAYER MET4 ;
    ANTENNAPARTIALMETALAREA 70.5 LAYER MET3 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA2 ;
    ANTENNAPARTIALCUTAREA 1.6929 LAYER VIA4 ;
    PORT
      LAYER MET5 ;
        RECT 0 78.5 65 89.5 ;
        RECT 0 3.788 1.5 15.212 ;
        RECT 0 3.753 1.476 15.247 ;
        RECT 0 3.707 1.43 15.293 ;
        RECT 0 3.661 1.384 15.339 ;
        RECT 0 3.615 1.338 15.385 ;
        RECT 0 3.569 1.292 15.431 ;
        RECT 0 3.523 1.246 15.477 ;
        RECT 0 3.5 1.2 15.5 ;
        RECT 0 17.288 1.5 28.712 ;
        RECT 0 17.253 1.476 28.747 ;
        RECT 0 17.207 1.43 28.793 ;
        RECT 0 17.161 1.384 28.839 ;
        RECT 0 17.115 1.338 28.885 ;
        RECT 0 17.069 1.292 28.931 ;
        RECT 0 17.023 1.246 28.977 ;
        RECT 0 17 1.2 29 ;
      LAYER MET4 ;
        RECT 0 79.483 6.5 88.517 ;
        RECT 0 79.443 6.466 88.557 ;
        RECT 0 79.397 6.42 88.603 ;
        RECT 0 79.351 6.374 88.649 ;
        RECT 0 79.305 6.328 88.695 ;
        RECT 0 79.259 6.282 88.741 ;
        RECT 0 79.213 6.236 88.787 ;
        RECT 0 79.167 6.19 88.833 ;
        RECT 0 79.121 6.144 88.879 ;
        RECT 0 79.075 6.098 88.925 ;
        RECT 0 79.029 6.052 88.971 ;
        RECT 0 78.983 6.006 89.017 ;
        RECT 0 78.937 5.96 89.063 ;
        RECT 0 78.891 5.914 89.109 ;
        RECT 0 78.845 5.868 89.155 ;
        RECT 0 78.799 5.822 89.201 ;
        RECT 0 78.753 5.776 89.247 ;
        RECT 0 78.707 5.73 89.293 ;
        RECT 0 78.661 5.684 89.339 ;
        RECT 0 78.615 5.638 89.385 ;
        RECT 0 78.569 5.592 89.431 ;
        RECT 0 78.523 5.546 89.477 ;
        RECT 0 78.5 5.5 89.5 ;
        RECT 0 3.788 1.5 15.212 ;
        RECT 0 3.753 1.476 15.247 ;
        RECT 0 3.707 1.43 15.293 ;
        RECT 0 3.661 1.384 15.339 ;
        RECT 0 3.615 1.338 15.385 ;
        RECT 0 3.569 1.292 15.431 ;
        RECT 0 3.523 1.246 15.477 ;
        RECT 0 3.5 1.2 15.5 ;
        RECT 0 17.288 1.5 28.712 ;
        RECT 0 17.253 1.476 28.747 ;
        RECT 0 17.207 1.43 28.793 ;
        RECT 0 17.161 1.384 28.839 ;
        RECT 0 17.115 1.338 28.885 ;
        RECT 0 17.069 1.292 28.931 ;
        RECT 0 17.023 1.246 28.977 ;
        RECT 0 17 1.2 29 ;
      LAYER MET3 ;
        RECT 0 79.483 6.5 88.517 ;
        RECT 0 79.443 6.466 88.557 ;
        RECT 0 79.397 6.42 88.603 ;
        RECT 0 79.351 6.374 88.649 ;
        RECT 0 79.305 6.328 88.695 ;
        RECT 0 79.259 6.282 88.741 ;
        RECT 0 79.213 6.236 88.787 ;
        RECT 0 79.167 6.19 88.833 ;
        RECT 0 79.121 6.144 88.879 ;
        RECT 0 79.075 6.098 88.925 ;
        RECT 0 79.029 6.052 88.971 ;
        RECT 0 78.983 6.006 89.017 ;
        RECT 0 78.937 5.96 89.063 ;
        RECT 0 78.891 5.914 89.109 ;
        RECT 0 78.845 5.868 89.155 ;
        RECT 0 78.799 5.822 89.201 ;
        RECT 0 78.753 5.776 89.247 ;
        RECT 0 78.707 5.73 89.293 ;
        RECT 0 78.661 5.684 89.339 ;
        RECT 0 78.615 5.638 89.385 ;
        RECT 0 78.569 5.592 89.431 ;
        RECT 0 78.523 5.546 89.477 ;
        RECT 0 78.5 5.5 89.5 ;
        RECT 0 3.788 1.5 15.212 ;
        RECT 0 3.753 1.476 15.247 ;
        RECT 0 3.707 1.43 15.293 ;
        RECT 0 3.661 1.384 15.339 ;
        RECT 0 3.615 1.338 15.385 ;
        RECT 0 3.569 1.292 15.431 ;
        RECT 0 3.523 1.246 15.477 ;
        RECT 0 3.5 1.2 15.5 ;
        RECT 0 17.288 1.5 28.712 ;
        RECT 0 17.253 1.476 28.747 ;
        RECT 0 17.207 1.43 28.793 ;
        RECT 0 17.161 1.384 28.839 ;
        RECT 0 17.115 1.338 28.885 ;
        RECT 0 17.069 1.292 28.931 ;
        RECT 0 17.023 1.246 28.977 ;
        RECT 0 17 1.2 29 ;
      LAYER MET2 ;
        RECT 0 17 65 29 ;
        RECT 0 3.5 65 15.5 ;
        RECT 59.805 3.5 60.995 29 ;
        RECT 54.225 3.5 55.415 29 ;
        RECT 48.645 3.5 49.835 29 ;
        RECT 43.065 3.5 44.255 29 ;
        RECT 37.485 3.5 38.675 29 ;
        RECT 31.905 3.5 33.095 29 ;
        RECT 26.325 3.5 27.515 29 ;
        RECT 20.745 3.5 21.935 29 ;
        RECT 15.165 3.5 16.355 29 ;
        RECT 9.585 3.5 10.775 29 ;
        RECT 4.005 3.5 5.195 29 ;
        RECT 0 78.5 65 89.5 ;
    END
  END VSSA
  OBS
    LAYER MET1 SPACING 0.09 ;
      RECT 0 -20 65 110 ;
    LAYER MET2 SPACING 0.1 ;
      RECT 57.175 107.675 65 110 ;
      RECT 0 107.675 7.825 110 ;
      RECT 0 107.675 65 108.825 ;
      RECT 0 -20 65 3.325 ;
      RECT 61.17 15.675 65 16.825 ;
      RECT 0 29.175 65 30.325 ;
      RECT 59.38 42.675 65 43.825 ;
      RECT 59.38 56.175 65 57.325 ;
      RECT 0 63.675 65 68.325 ;
      RECT 0 77.175 65 78.325 ;
      RECT 0 89.675 65 90.825 ;
      RECT 0 98.175 65 99.325 ;
      RECT 55.59 15.675 59.63 16.825 ;
      RECT 53.8 42.675 55.84 43.825 ;
      RECT 53.8 56.175 55.84 57.325 ;
      RECT 50.01 15.675 54.05 16.825 ;
      RECT 48.22 42.675 50.26 43.825 ;
      RECT 48.22 56.175 50.26 57.325 ;
      RECT 44.43 15.675 48.47 16.825 ;
      RECT 42.64 42.675 44.68 43.825 ;
      RECT 42.64 56.175 44.68 57.325 ;
      RECT 38.85 15.675 42.89 16.825 ;
      RECT 37.06 42.675 39.1 43.825 ;
      RECT 37.06 56.175 39.1 57.325 ;
      RECT 33.27 15.675 37.31 16.825 ;
      RECT 31.48 42.675 33.52 43.825 ;
      RECT 31.48 56.175 33.52 57.325 ;
      RECT 27.69 15.675 31.73 16.825 ;
      RECT 25.9 42.675 27.94 43.825 ;
      RECT 25.9 56.175 27.94 57.325 ;
      RECT 22.11 15.675 26.15 16.825 ;
      RECT 20.32 42.675 22.36 43.825 ;
      RECT 20.32 56.175 22.36 57.325 ;
      RECT 16.53 15.675 20.57 16.825 ;
      RECT 14.74 42.675 16.78 43.825 ;
      RECT 14.74 56.175 16.78 57.325 ;
      RECT 10.95 15.675 14.99 16.825 ;
      RECT 9.16 42.675 11.2 43.825 ;
      RECT 9.16 56.175 11.2 57.325 ;
      RECT 5.37 15.675 9.41 16.825 ;
      RECT 0 42.675 5.62 43.825 ;
      RECT 0 56.175 5.62 57.325 ;
      RECT 0 15.675 3.83 16.825 ;
    LAYER MET3 SPACING 0.1 ;
      RECT 61.175 -20 65 3.335 ;
      RECT 1.375 -20 3.825 3.335 ;
      RECT 0 -20 3.825 3.325 ;
      RECT 0 -20 65 -0.175 ;
      RECT 63.8 3.5 65 15.5 ;
      RECT 63.776 3.512 65 15.488 ;
      RECT 63.73 3.547 65 15.453 ;
      RECT 63.684 3.593 65 15.407 ;
      RECT 63.638 3.639 65 15.361 ;
      RECT 63.592 3.685 65 15.315 ;
      RECT 63.546 3.731 65 15.269 ;
      RECT 63.5 3.777 65 15.223 ;
      RECT 63.8 17 65 29 ;
      RECT 63.776 17.012 65 28.988 ;
      RECT 63.73 17.047 65 28.953 ;
      RECT 63.684 17.093 65 28.907 ;
      RECT 63.638 17.139 65 28.861 ;
      RECT 63.592 17.185 65 28.815 ;
      RECT 63.546 17.231 65 28.769 ;
      RECT 63.5 17.277 65 28.723 ;
      RECT 63.8 30.5 65 42.5 ;
      RECT 63.776 30.512 65 42.488 ;
      RECT 63.73 30.547 65 42.453 ;
      RECT 63.684 30.593 65 42.407 ;
      RECT 63.638 30.639 65 42.361 ;
      RECT 63.592 30.685 65 42.315 ;
      RECT 63.546 30.731 65 42.269 ;
      RECT 63.5 30.777 65 42.223 ;
      RECT 63.8 44 65 56 ;
      RECT 63.776 44.012 65 55.988 ;
      RECT 63.73 44.047 65 55.953 ;
      RECT 63.684 44.093 65 55.907 ;
      RECT 63.638 44.139 65 55.861 ;
      RECT 63.592 44.185 65 55.815 ;
      RECT 63.546 44.231 65 55.769 ;
      RECT 63.5 44.277 65 55.723 ;
      RECT 63.8 57.5 65 63.5 ;
      RECT 63.776 57.512 65 63.488 ;
      RECT 63.73 57.547 65 63.453 ;
      RECT 63.684 57.593 65 63.407 ;
      RECT 63.638 57.639 65 63.361 ;
      RECT 63.592 57.685 65 63.315 ;
      RECT 63.546 57.731 65 63.269 ;
      RECT 63.5 57.777 65 63.223 ;
      RECT 62.175 63.665 65 68.335 ;
      RECT 57.175 63.675 65 68.325 ;
      RECT 63.8 68.5 65 77 ;
      RECT 63.776 68.512 65 76.988 ;
      RECT 63.73 68.547 65 76.953 ;
      RECT 63.684 68.593 65 76.907 ;
      RECT 63.638 68.639 65 76.861 ;
      RECT 63.592 68.685 65 76.815 ;
      RECT 63.546 68.731 65 76.769 ;
      RECT 63.5 68.777 65 76.723 ;
      RECT 57.175 77.175 65 78.335 ;
      RECT 62.175 77.165 65 78.335 ;
      RECT 59.466 78.517 59.5 89.483 ;
      RECT 59.42 78.557 59.466 89.443 ;
      RECT 59.374 78.603 59.42 89.397 ;
      RECT 59.328 78.649 59.374 89.351 ;
      RECT 59.282 78.695 59.328 89.305 ;
      RECT 59.236 78.741 59.282 89.259 ;
      RECT 59.19 78.787 59.236 89.213 ;
      RECT 59.144 78.833 59.19 89.167 ;
      RECT 59.098 78.879 59.144 89.121 ;
      RECT 59.052 78.925 59.098 89.075 ;
      RECT 59.006 78.971 59.052 89.029 ;
      RECT 58.96 79.017 59.006 88.983 ;
      RECT 58.914 79.063 58.96 88.937 ;
      RECT 58.868 79.109 58.914 88.891 ;
      RECT 58.822 79.155 58.868 88.845 ;
      RECT 58.776 79.201 58.822 88.799 ;
      RECT 58.73 79.247 58.776 88.753 ;
      RECT 58.684 79.293 58.73 88.707 ;
      RECT 58.638 79.339 58.684 88.661 ;
      RECT 58.592 79.385 58.638 88.615 ;
      RECT 58.546 79.431 58.592 88.569 ;
      RECT 58.5 79.477 58.546 88.523 ;
      RECT 59.5 78.5 65 89.5 ;
      RECT 59.466 91.017 59.5 97.983 ;
      RECT 59.42 91.057 59.466 97.943 ;
      RECT 59.374 91.103 59.42 97.897 ;
      RECT 59.328 91.149 59.374 97.851 ;
      RECT 59.282 91.195 59.328 97.805 ;
      RECT 59.236 91.241 59.282 97.759 ;
      RECT 59.19 91.287 59.236 97.713 ;
      RECT 59.144 91.333 59.19 97.667 ;
      RECT 59.098 91.379 59.144 97.621 ;
      RECT 59.052 91.425 59.098 97.575 ;
      RECT 59.006 91.471 59.052 97.529 ;
      RECT 58.96 91.517 59.006 97.483 ;
      RECT 58.914 91.563 58.96 97.437 ;
      RECT 58.868 91.609 58.914 97.391 ;
      RECT 58.822 91.655 58.868 97.345 ;
      RECT 58.776 91.701 58.822 97.299 ;
      RECT 58.73 91.747 58.776 97.253 ;
      RECT 58.684 91.793 58.73 97.207 ;
      RECT 58.638 91.839 58.684 97.161 ;
      RECT 58.592 91.885 58.638 97.115 ;
      RECT 58.546 91.931 58.592 97.069 ;
      RECT 58.5 91.977 58.546 97.023 ;
      RECT 59.5 91 65 98 ;
      RECT 59.466 99.517 59.5 107.483 ;
      RECT 59.42 99.557 59.466 107.443 ;
      RECT 59.374 99.603 59.42 107.397 ;
      RECT 59.328 99.649 59.374 107.351 ;
      RECT 59.282 99.695 59.328 107.305 ;
      RECT 59.236 99.741 59.282 107.259 ;
      RECT 59.19 99.787 59.236 107.213 ;
      RECT 59.144 99.833 59.19 107.167 ;
      RECT 59.098 99.879 59.144 107.121 ;
      RECT 59.052 99.925 59.098 107.075 ;
      RECT 59.006 99.971 59.052 107.029 ;
      RECT 58.96 100.017 59.006 106.983 ;
      RECT 58.914 100.063 58.96 106.937 ;
      RECT 58.868 100.109 58.914 106.891 ;
      RECT 58.822 100.155 58.868 106.845 ;
      RECT 58.776 100.201 58.822 106.799 ;
      RECT 58.73 100.247 58.776 106.753 ;
      RECT 58.684 100.293 58.73 106.707 ;
      RECT 58.638 100.339 58.684 106.661 ;
      RECT 58.592 100.385 58.638 106.615 ;
      RECT 58.546 100.431 58.592 106.569 ;
      RECT 58.5 100.477 58.546 106.523 ;
      RECT 59.5 99.5 65 107.5 ;
      RECT 1.375 63.665 2.825 68.335 ;
      RECT 0 63.675 7.825 68.325 ;
      RECT 5.675 77.175 7.825 78.335 ;
      RECT 0 77.175 7.825 78.325 ;
      RECT 1.375 77.165 2.825 78.325 ;
      RECT 5.675 89.665 7.825 90.835 ;
      RECT 0 89.675 7.825 90.825 ;
      RECT 5.675 98.165 7.825 99.335 ;
      RECT 0 98.175 7.825 99.325 ;
      RECT 0 107.675 7.825 110 ;
      RECT 5.675 107.665 7.825 110 ;
      RECT 1.375 15.665 2.825 16.835 ;
      RECT 0 15.675 2.825 16.825 ;
      RECT 1.375 29.165 2.825 30.335 ;
      RECT 0 29.175 2.825 30.325 ;
      RECT 1.375 42.665 2.825 43.835 ;
      RECT 0 42.675 2.825 43.825 ;
      RECT 1.375 56.165 2.825 57.335 ;
      RECT 0 56.175 2.825 57.325 ;
      RECT 62.175 15.665 65 16.835 ;
      RECT 62.175 29.165 65 30.335 ;
      RECT 62.175 42.665 65 43.835 ;
      RECT 62.175 56.165 65 57.335 ;
      RECT 57.175 89.665 65 90.835 ;
      RECT 57.175 98.165 65 99.335 ;
      RECT 57.175 107.665 65 110 ;
      RECT 50.675 29.165 56.825 29.325 ;
      RECT 53.79 42.665 55.85 43.325 ;
      RECT 53.79 56.165 55.85 57.325 ;
      RECT 44.515 63.675 45.825 68.325 ;
      RECT 44.515 77.175 45.825 78.335 ;
      RECT 44.515 89.665 45.825 90.835 ;
      RECT 44.515 98.165 45.825 99.335 ;
      RECT 44.515 107.665 45.825 108.825 ;
      RECT 36.675 29.165 42.825 29.325 ;
      RECT 42.63 42.665 42.825 43.325 ;
      RECT 42.63 56.165 42.825 57.325 ;
      RECT 37.05 42.665 39.11 43.325 ;
      RECT 37.05 56.165 39.11 57.325 ;
      RECT 31.835 63.675 33.095 68.325 ;
      RECT 31.835 77.175 33.095 78.335 ;
      RECT 31.835 89.665 33.095 90.835 ;
      RECT 31.835 98.165 33.095 99.335 ;
      RECT 31.835 107.665 33.095 108.825 ;
      RECT 22.675 29.165 28.825 29.325 ;
      RECT 25.89 42.665 27.95 43.325 ;
      RECT 25.89 56.165 27.95 57.325 ;
      RECT 19.175 63.675 20.485 68.325 ;
      RECT 19.175 77.175 20.485 78.335 ;
      RECT 19.175 89.665 20.485 90.835 ;
      RECT 19.175 98.165 20.485 99.335 ;
      RECT 19.175 107.665 20.485 108.825 ;
      RECT 8.675 29.165 14.825 29.325 ;
      RECT 9.15 42.665 11.21 43.325 ;
      RECT 9.15 56.165 11.21 57.325 ;
    LAYER MET4 SPACING 0.1 ;
      RECT 57.175 77.175 65 110 ;
      RECT 62.175 -20 65 110 ;
      RECT 0 107.675 7.825 110 ;
      RECT 6.675 77.175 7.825 110 ;
      RECT 5.675 107.652 7.825 110 ;
      RECT 6.641 106.692 7.825 110 ;
      RECT 5.721 107.606 7.825 110 ;
      RECT 6.595 106.732 7.825 110 ;
      RECT 5.767 107.56 7.825 110 ;
      RECT 6.549 106.778 7.825 110 ;
      RECT 5.813 107.514 7.825 110 ;
      RECT 6.503 106.824 7.825 110 ;
      RECT 5.859 107.468 7.825 110 ;
      RECT 6.457 106.87 7.825 110 ;
      RECT 5.905 107.422 7.825 110 ;
      RECT 6.411 106.916 7.825 110 ;
      RECT 5.951 107.376 7.825 110 ;
      RECT 6.365 106.962 7.825 110 ;
      RECT 5.997 107.33 7.825 110 ;
      RECT 6.319 107.008 7.825 110 ;
      RECT 6.043 107.284 7.825 110 ;
      RECT 6.273 107.054 7.825 110 ;
      RECT 6.089 107.238 7.825 110 ;
      RECT 6.227 107.1 7.825 110 ;
      RECT 6.135 107.192 7.825 110 ;
      RECT 6.181 107.146 7.825 110 ;
      RECT 6.641 97.192 7.825 100.308 ;
      RECT 6.595 97.232 7.825 100.268 ;
      RECT 6.549 97.278 7.825 100.222 ;
      RECT 6.503 97.324 7.825 100.176 ;
      RECT 6.457 97.37 7.825 100.13 ;
      RECT 6.411 97.416 7.825 100.084 ;
      RECT 6.365 97.462 7.825 100.038 ;
      RECT 6.319 97.508 7.825 99.992 ;
      RECT 6.273 97.554 7.825 99.946 ;
      RECT 6.227 97.6 7.825 99.9 ;
      RECT 6.181 97.646 7.825 99.854 ;
      RECT 6.135 97.692 7.825 99.808 ;
      RECT 6.089 97.738 7.825 99.762 ;
      RECT 6.043 97.784 7.825 99.716 ;
      RECT 5.997 97.83 7.825 99.67 ;
      RECT 5.951 97.876 7.825 99.624 ;
      RECT 5.905 97.922 7.825 99.578 ;
      RECT 5.859 97.968 7.825 99.532 ;
      RECT 5.813 98.014 7.825 99.486 ;
      RECT 5.767 98.06 7.825 99.44 ;
      RECT 5.721 98.106 7.825 99.394 ;
      RECT 5.675 98.152 7.825 99.348 ;
      RECT 0 98.175 7.825 99.325 ;
      RECT 6.641 88.692 7.825 91.808 ;
      RECT 6.595 88.732 7.825 91.768 ;
      RECT 6.549 88.778 7.825 91.722 ;
      RECT 6.503 88.824 7.825 91.676 ;
      RECT 6.457 88.87 7.825 91.63 ;
      RECT 6.411 88.916 7.825 91.584 ;
      RECT 6.365 88.962 7.825 91.538 ;
      RECT 6.319 89.008 7.825 91.492 ;
      RECT 6.273 89.054 7.825 91.446 ;
      RECT 6.227 89.1 7.825 91.4 ;
      RECT 6.181 89.146 7.825 91.354 ;
      RECT 6.135 89.192 7.825 91.308 ;
      RECT 6.089 89.238 7.825 91.262 ;
      RECT 6.043 89.284 7.825 91.216 ;
      RECT 5.997 89.33 7.825 91.17 ;
      RECT 5.951 89.376 7.825 91.124 ;
      RECT 5.905 89.422 7.825 91.078 ;
      RECT 5.859 89.468 7.825 91.032 ;
      RECT 5.813 89.514 7.825 90.986 ;
      RECT 5.767 89.56 7.825 90.94 ;
      RECT 5.721 89.606 7.825 90.894 ;
      RECT 5.675 89.652 7.825 90.848 ;
      RECT 0 89.675 7.825 90.825 ;
      RECT 6.641 77.175 7.825 79.308 ;
      RECT 6.595 77.175 7.825 79.268 ;
      RECT 6.549 77.175 7.825 79.222 ;
      RECT 6.503 77.175 7.825 79.176 ;
      RECT 6.457 77.175 7.825 79.13 ;
      RECT 6.411 77.175 7.825 79.084 ;
      RECT 6.365 77.175 7.825 79.038 ;
      RECT 6.319 77.175 7.825 78.992 ;
      RECT 6.273 77.175 7.825 78.946 ;
      RECT 6.227 77.175 7.825 78.9 ;
      RECT 6.181 77.175 7.825 78.854 ;
      RECT 6.135 77.175 7.825 78.808 ;
      RECT 6.089 77.175 7.825 78.762 ;
      RECT 6.043 77.175 7.825 78.716 ;
      RECT 5.997 77.175 7.825 78.67 ;
      RECT 5.951 77.175 7.825 78.624 ;
      RECT 5.905 77.175 7.825 78.578 ;
      RECT 5.859 77.175 7.825 78.532 ;
      RECT 5.813 77.175 7.825 78.486 ;
      RECT 5.767 77.175 7.825 78.44 ;
      RECT 5.721 77.175 7.825 78.394 ;
      RECT 5.675 77.175 7.825 78.348 ;
      RECT 0 77.175 7.825 78.325 ;
      RECT 1.375 77.152 2.825 78.325 ;
      RECT 1.675 -20 2.825 78.325 ;
      RECT 1.421 77.106 2.825 78.325 ;
      RECT 1.651 76.887 2.825 78.325 ;
      RECT 1.467 77.06 2.825 78.325 ;
      RECT 1.605 76.922 2.825 78.325 ;
      RECT 1.513 77.014 2.825 78.325 ;
      RECT 1.559 76.968 2.825 78.325 ;
      RECT 1.651 63.387 2.825 68.613 ;
      RECT 1.605 63.422 2.825 68.578 ;
      RECT 1.559 63.468 2.825 68.532 ;
      RECT 1.513 63.514 2.825 68.486 ;
      RECT 1.467 63.56 2.825 68.44 ;
      RECT 1.421 63.606 2.825 68.394 ;
      RECT 1.375 63.652 2.825 68.348 ;
      RECT 57.175 63.675 65 68.325 ;
      RECT 0 63.675 7.825 68.325 ;
      RECT 1.651 55.887 2.825 57.613 ;
      RECT 1.605 55.922 2.825 57.578 ;
      RECT 1.559 55.968 2.825 57.532 ;
      RECT 1.513 56.014 2.825 57.486 ;
      RECT 1.467 56.06 2.825 57.44 ;
      RECT 1.421 56.106 2.825 57.394 ;
      RECT 1.375 56.152 2.825 57.348 ;
      RECT 0 56.175 2.825 57.325 ;
      RECT 1.651 42.387 2.825 44.113 ;
      RECT 1.605 42.422 2.825 44.078 ;
      RECT 1.559 42.468 2.825 44.032 ;
      RECT 1.513 42.514 2.825 43.986 ;
      RECT 1.467 42.56 2.825 43.94 ;
      RECT 1.421 42.606 2.825 43.894 ;
      RECT 1.375 42.652 2.825 43.848 ;
      RECT 0 42.675 2.825 43.825 ;
      RECT 1.651 28.887 2.825 30.613 ;
      RECT 1.605 28.922 2.825 30.578 ;
      RECT 1.559 28.968 2.825 30.532 ;
      RECT 1.513 29.014 2.825 30.486 ;
      RECT 1.467 29.06 2.825 30.44 ;
      RECT 1.421 29.106 2.825 30.394 ;
      RECT 1.375 29.152 2.825 30.348 ;
      RECT 0 29.175 2.825 30.325 ;
      RECT 1.651 15.387 2.825 17.113 ;
      RECT 1.605 15.422 2.825 17.078 ;
      RECT 1.559 15.468 2.825 17.032 ;
      RECT 1.513 15.514 2.825 16.986 ;
      RECT 1.467 15.56 2.825 16.94 ;
      RECT 1.421 15.606 2.825 16.894 ;
      RECT 1.375 15.652 2.825 16.848 ;
      RECT 0 15.675 2.825 16.825 ;
      RECT 62.141 -20 65 4.308 ;
      RECT 1.675 -20 2.871 4.302 ;
      RECT 62.095 -20 65 4.268 ;
      RECT 1.675 -20 2.917 4.256 ;
      RECT 62.049 -20 65 4.222 ;
      RECT 1.675 -20 2.963 4.21 ;
      RECT 62.003 -20 65 4.176 ;
      RECT 1.675 -20 3.009 4.164 ;
      RECT 61.957 -20 65 4.13 ;
      RECT 1.675 -20 3.055 4.118 ;
      RECT 61.911 -20 65 4.084 ;
      RECT 1.675 -20 3.101 4.072 ;
      RECT 61.865 -20 65 4.038 ;
      RECT 1.675 -20 3.147 4.026 ;
      RECT 61.819 -20 65 3.992 ;
      RECT 1.675 -20 3.193 3.98 ;
      RECT 61.773 -20 65 3.946 ;
      RECT 1.675 -20 3.239 3.934 ;
      RECT 61.727 -20 65 3.9 ;
      RECT 1.675 -20 3.285 3.888 ;
      RECT 61.681 -20 65 3.854 ;
      RECT 1.675 -20 3.331 3.842 ;
      RECT 61.635 -20 65 3.808 ;
      RECT 1.675 -20 3.377 3.796 ;
      RECT 61.589 -20 65 3.762 ;
      RECT 1.675 -20 3.423 3.75 ;
      RECT 61.543 -20 65 3.716 ;
      RECT 1.675 -20 3.469 3.704 ;
      RECT 61.497 -20 65 3.67 ;
      RECT 1.675 -20 3.515 3.658 ;
      RECT 61.451 -20 65 3.624 ;
      RECT 1.651 -20 3.515 3.613 ;
      RECT 1.651 -20 3.561 3.612 ;
      RECT 61.405 -20 65 3.578 ;
      RECT 1.605 -20 3.561 3.578 ;
      RECT 1.605 -20 3.607 3.566 ;
      RECT 61.359 -20 65 3.532 ;
      RECT 1.559 -20 3.607 3.532 ;
      RECT 1.559 -20 3.653 3.52 ;
      RECT 61.313 -20 65 3.486 ;
      RECT 1.513 -20 3.653 3.486 ;
      RECT 1.513 -20 3.699 3.474 ;
      RECT 61.267 -20 65 3.44 ;
      RECT 1.467 -20 3.699 3.44 ;
      RECT 1.467 -20 3.745 3.428 ;
      RECT 61.221 -20 65 3.394 ;
      RECT 1.421 -20 3.745 3.394 ;
      RECT 1.421 -20 3.791 3.382 ;
      RECT 61.175 -20 65 3.348 ;
      RECT 1.375 -20 3.791 3.348 ;
      RECT 1.375 -20 3.825 3.342 ;
      RECT 0 -20 3.825 3.325 ;
      RECT 0 -20 65 -0.175 ;
      RECT 50.675 9.175 56.825 15.325 ;
      RECT 50.675 23.175 56.825 29.325 ;
      RECT 50.675 37.175 56.825 43.325 ;
      RECT 50.675 51.175 56.825 57.325 ;
      RECT 44.515 63.675 45.825 68.325 ;
      RECT 44.515 77.175 45.825 108.825 ;
      RECT 36.675 9.175 42.825 15.325 ;
      RECT 36.675 23.175 42.825 29.325 ;
      RECT 36.675 37.175 42.825 43.325 ;
      RECT 36.675 51.175 42.825 57.325 ;
      RECT 31.835 63.675 33.095 68.325 ;
      RECT 31.835 77.175 33.095 108.825 ;
      RECT 22.675 9.175 28.825 15.325 ;
      RECT 22.675 23.175 28.825 29.325 ;
      RECT 22.675 37.175 28.825 43.325 ;
      RECT 22.675 51.175 28.825 57.325 ;
      RECT 19.175 63.675 20.485 68.325 ;
      RECT 19.175 77.175 20.485 108.825 ;
      RECT 8.675 9.175 14.825 15.325 ;
      RECT 8.675 23.175 14.825 29.325 ;
      RECT 8.675 37.175 14.825 43.325 ;
      RECT 8.675 51.175 14.825 57.325 ;
    LAYER MET5 SPACING 0.1 ;
      RECT 57.165 77.165 65 78.17 ;
      RECT 62.165 -20 65 78.17 ;
      RECT 0 77.33 7.835 78.17 ;
      RECT 1.714 77.165 7.835 78.17 ;
      RECT 1.53 77.307 7.835 78.17 ;
      RECT 1.668 77.169 7.835 78.17 ;
      RECT 1.576 77.261 7.835 78.17 ;
      RECT 1.622 77.215 7.835 78.17 ;
      RECT 1.714 77.123 2.835 78.17 ;
      RECT 1.83 -20 2.835 78.17 ;
      RECT 1.76 77.077 2.835 78.17 ;
      RECT 1.806 77.042 2.835 78.17 ;
      RECT 1.806 63.542 2.835 68.458 ;
      RECT 1.76 63.577 2.835 68.423 ;
      RECT 1.714 63.623 2.835 68.377 ;
      RECT 57.165 63.665 65 68.335 ;
      RECT 1.714 63.665 7.835 68.335 ;
      RECT 1.668 63.669 7.835 68.331 ;
      RECT 1.622 63.715 7.835 68.285 ;
      RECT 1.576 63.761 7.835 68.239 ;
      RECT 1.53 63.807 7.835 68.193 ;
      RECT 0 63.83 7.835 68.17 ;
      RECT 1.806 56.042 2.835 57.458 ;
      RECT 1.76 56.077 2.835 57.423 ;
      RECT 1.714 56.123 2.835 57.377 ;
      RECT 1.668 56.169 2.835 57.331 ;
      RECT 1.622 56.215 2.835 57.285 ;
      RECT 1.576 56.261 2.835 57.239 ;
      RECT 1.53 56.307 2.835 57.193 ;
      RECT 0 56.33 2.835 57.17 ;
      RECT 1.806 42.542 2.835 43.958 ;
      RECT 1.76 42.577 2.835 43.923 ;
      RECT 1.714 42.623 2.835 43.877 ;
      RECT 1.668 42.669 2.835 43.831 ;
      RECT 1.622 42.715 2.835 43.785 ;
      RECT 1.576 42.761 2.835 43.739 ;
      RECT 1.53 42.807 2.835 43.693 ;
      RECT 0 42.83 2.835 43.67 ;
      RECT 1.806 29.042 2.835 30.458 ;
      RECT 1.76 29.077 2.835 30.423 ;
      RECT 1.714 29.123 2.835 30.377 ;
      RECT 1.668 29.169 2.835 30.331 ;
      RECT 1.622 29.215 2.835 30.285 ;
      RECT 1.576 29.261 2.835 30.239 ;
      RECT 1.53 29.307 2.835 30.193 ;
      RECT 0 29.33 2.835 30.17 ;
      RECT 1.806 15.542 2.835 16.958 ;
      RECT 1.76 15.577 2.835 16.923 ;
      RECT 1.714 15.623 2.835 16.877 ;
      RECT 1.668 15.669 2.835 16.831 ;
      RECT 1.622 15.715 2.835 16.785 ;
      RECT 1.576 15.761 2.835 16.739 ;
      RECT 1.53 15.807 2.835 16.693 ;
      RECT 0 15.83 2.835 16.67 ;
      RECT 62.131 -20 65 4.318 ;
      RECT 1.83 -20 2.881 4.312 ;
      RECT 62.085 -20 65 4.278 ;
      RECT 1.83 -20 2.927 4.266 ;
      RECT 62.039 -20 65 4.232 ;
      RECT 1.83 -20 2.973 4.22 ;
      RECT 61.993 -20 65 4.186 ;
      RECT 1.83 -20 3.019 4.174 ;
      RECT 61.947 -20 65 4.14 ;
      RECT 1.83 -20 3.065 4.128 ;
      RECT 61.901 -20 65 4.094 ;
      RECT 1.83 -20 3.111 4.082 ;
      RECT 61.855 -20 65 4.048 ;
      RECT 1.83 -20 3.157 4.036 ;
      RECT 61.809 -20 65 4.002 ;
      RECT 1.83 -20 3.203 3.99 ;
      RECT 61.763 -20 65 3.956 ;
      RECT 1.83 -20 3.249 3.944 ;
      RECT 61.717 -20 65 3.91 ;
      RECT 1.83 -20 3.295 3.898 ;
      RECT 61.671 -20 65 3.864 ;
      RECT 1.83 -20 3.341 3.852 ;
      RECT 61.625 -20 65 3.818 ;
      RECT 1.83 -20 3.387 3.806 ;
      RECT 61.579 -20 65 3.772 ;
      RECT 1.83 -20 3.433 3.76 ;
      RECT 61.533 -20 65 3.726 ;
      RECT 1.83 -20 3.479 3.714 ;
      RECT 61.487 -20 65 3.68 ;
      RECT 1.83 -20 3.525 3.668 ;
      RECT 61.441 -20 65 3.634 ;
      RECT 1.83 -20 3.571 3.622 ;
      RECT 61.395 -20 65 3.588 ;
      RECT 1.83 -20 3.617 3.576 ;
      RECT 61.349 -20 65 3.542 ;
      RECT 1.83 -20 3.663 3.53 ;
      RECT 61.303 -20 65 3.496 ;
      RECT 1.83 -20 3.709 3.484 ;
      RECT 1.806 -20 3.709 3.458 ;
      RECT 61.257 -20 65 3.45 ;
      RECT 1.806 -20 3.755 3.438 ;
      RECT 1.76 -20 3.755 3.423 ;
      RECT 61.211 -20 65 3.404 ;
      RECT 1.76 -20 3.801 3.392 ;
      RECT 1.714 -20 3.801 3.377 ;
      RECT 61.165 -20 65 3.358 ;
      RECT 1.714 -20 3.835 3.352 ;
      RECT 1.668 -20 3.835 3.331 ;
      RECT 1.622 -20 3.835 3.285 ;
      RECT 1.576 -20 3.835 3.239 ;
      RECT 1.53 -20 3.835 3.193 ;
      RECT 0 -20 3.835 3.17 ;
      RECT 0 -20 65 -0.165 ;
      RECT 57.33 107.83 65 110 ;
      RECT 57.165 107.83 65 108.67 ;
      RECT 3 68.5 62 77 ;
      RECT 8 0 57 77 ;
      RECT 4 0 61 63.5 ;
      RECT 61.966 4.483 62 63.5 ;
      RECT 61.92 4.443 61.966 63.5 ;
      RECT 61.874 4.397 61.92 63.5 ;
      RECT 61.828 4.351 61.874 63.5 ;
      RECT 61.782 4.305 61.828 63.5 ;
      RECT 61.736 4.259 61.782 63.5 ;
      RECT 61.69 4.213 61.736 63.5 ;
      RECT 61.644 4.167 61.69 63.5 ;
      RECT 61.598 4.121 61.644 63.5 ;
      RECT 61.552 4.075 61.598 63.5 ;
      RECT 61.506 4.029 61.552 63.5 ;
      RECT 61.46 3.983 61.506 63.5 ;
      RECT 61.414 3.937 61.46 63.5 ;
      RECT 61.368 3.891 61.414 63.5 ;
      RECT 61.322 3.845 61.368 63.5 ;
      RECT 61.276 3.799 61.322 63.5 ;
      RECT 61.23 3.753 61.276 63.5 ;
      RECT 61.184 3.707 61.23 63.5 ;
      RECT 61.138 3.661 61.184 63.5 ;
      RECT 61.092 3.615 61.138 63.5 ;
      RECT 61.046 3.569 61.092 63.5 ;
      RECT 61 3.523 61.046 63.5 ;
      RECT 3.966 3.517 4 63.5 ;
      RECT 3.92 3.557 3.966 63.5 ;
      RECT 3.874 3.603 3.92 63.5 ;
      RECT 3.828 3.649 3.874 63.5 ;
      RECT 3.782 3.695 3.828 63.5 ;
      RECT 3.736 3.741 3.782 63.5 ;
      RECT 3.69 3.787 3.736 63.5 ;
      RECT 3.644 3.833 3.69 63.5 ;
      RECT 3.598 3.879 3.644 63.5 ;
      RECT 3.552 3.925 3.598 63.5 ;
      RECT 3.506 3.971 3.552 63.5 ;
      RECT 3.46 4.017 3.506 63.5 ;
      RECT 3.414 4.063 3.46 63.5 ;
      RECT 3.368 4.109 3.414 63.5 ;
      RECT 3.322 4.155 3.368 63.5 ;
      RECT 3.276 4.201 3.322 63.5 ;
      RECT 3.23 4.247 3.276 63.5 ;
      RECT 3.184 4.293 3.23 63.5 ;
      RECT 3.138 4.339 3.184 63.5 ;
      RECT 3.092 4.385 3.138 63.5 ;
      RECT 3.046 4.431 3.092 63.5 ;
      RECT 3 4.477 3.046 63.5 ;
      RECT 0 107.83 7.67 110 ;
      RECT 0 107.83 7.835 108.67 ;
      RECT 57.165 89.83 65 90.67 ;
      RECT 57.165 98.33 65 99.17 ;
      RECT 44.505 77.165 45.835 78.17 ;
      RECT 44.505 89.83 45.835 90.67 ;
      RECT 44.505 98.33 45.835 99.17 ;
      RECT 44.505 107.83 45.835 108.67 ;
      RECT 31.825 77.165 33.105 78.17 ;
      RECT 31.825 89.83 33.105 90.67 ;
      RECT 31.825 98.33 33.105 99.17 ;
      RECT 31.825 107.83 33.105 108.67 ;
      RECT 19.165 77.165 20.495 78.17 ;
      RECT 19.165 89.83 20.495 90.67 ;
      RECT 19.165 98.33 20.495 99.17 ;
      RECT 19.165 107.83 20.495 108.67 ;
      RECT 0 89.83 7.835 90.67 ;
      RECT 0 98.33 7.835 99.17 ;
    LAYER T4M2 SPACING 0.4 ;
      RECT 64.584 -20 65 0.307 ;
      RECT 0 -20 0.428 0.295 ;
      RECT 64.538 -20 65 0.261 ;
      RECT 0 -20 0.474 0.249 ;
      RECT 64.492 -20 65 0.215 ;
      RECT 0 -20 0.52 0.203 ;
      RECT 64.446 -20 65 0.169 ;
      RECT 0 -20 0.566 0.157 ;
      RECT 64.4 -20 65 0.123 ;
      RECT 0 -20 0.6 0.117 ;
      RECT 0 -20 65 -3.4 ;
      RECT 57.6 108.1 65 110 ;
      RECT 0 108.1 7.4 110 ;
    LAYER RDL SPACING 2 ;
      RECT 0 -20 65 -5 ;
      RECT 0 82 65 110 ;
      RECT 3 4.5 62 63.5 ;
  END
END P65_1233_VDD1A

MACRO P65_1233_VDD3
  CLASS PAD ;
  ORIGIN 0 20 ;
  FOREIGN P65_1233_VDD3 0 -20 ;
  SIZE 65 BY 130 ;
  SYMMETRY X Y R90 ;
  SITE IOSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER MET5 ;
        RECT 8 109 57 110 ;
      LAYER MET4 ;
        RECT 8 109 57 110 ;
      LAYER MET3 ;
        RECT 8 109 57 110 ;
      LAYER MET2 ;
        RECT 8 99.5 57 110 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 99.5 65 107.5 ;
      LAYER T4M2 ;
        RECT 57 4.532 61.9 65.968 ;
        RECT 57 4.497 61.875 66.003 ;
        RECT 57 4.451 61.829 66.049 ;
        RECT 57 4.405 61.783 66.095 ;
        RECT 57 4.359 61.737 66.141 ;
        RECT 57 4.313 61.691 66.187 ;
        RECT 57 4.267 61.645 66.233 ;
        RECT 57 4.221 61.599 66.279 ;
        RECT 57 4.175 61.553 66.325 ;
        RECT 57 4.129 61.507 66.371 ;
        RECT 57 4.083 61.461 66.417 ;
        RECT 57 4.037 61.415 66.463 ;
        RECT 57 3.991 61.369 66.509 ;
        RECT 57 3.945 61.323 66.555 ;
        RECT 57 3.899 61.277 66.601 ;
        RECT 57 3.853 61.231 66.647 ;
        RECT 57 3.807 61.185 66.693 ;
        RECT 57 3.761 61.139 66.739 ;
        RECT 57 3.715 61.093 66.785 ;
        RECT 57 3.669 61.047 66.831 ;
        RECT 57 3.623 61.001 66.877 ;
        RECT 4.045 57.5 60.955 66.9 ;
        RECT 57 3.595 60.955 66.9 ;
        RECT 4.045 3.577 60.946 9 ;
        RECT 57 3.568 60.946 66.9 ;
        RECT 4.091 3.549 60.9 9 ;
        RECT 3.1 43.5 61.9 51 ;
        RECT 3.1 29.5 61.9 37 ;
        RECT 3.1 15.5 61.9 23 ;
        RECT 4.1 0.1 60.9 9 ;
        RECT 43 0.1 50.5 66.9 ;
        RECT 29 0.1 36.5 66.9 ;
        RECT 15 0.1 22.5 66.9 ;
        RECT 3.1 4.522 8.5 65.978 ;
        RECT 4.02 3.612 8.5 66.888 ;
        RECT 3.974 3.648 8.5 66.852 ;
        RECT 3.928 3.694 8.5 66.806 ;
        RECT 3.882 3.74 8.5 66.76 ;
        RECT 3.836 3.786 8.5 66.714 ;
        RECT 3.79 3.832 8.5 66.668 ;
        RECT 3.744 3.878 8.5 66.622 ;
        RECT 3.698 3.924 8.5 66.576 ;
        RECT 3.652 3.97 8.5 66.53 ;
        RECT 3.606 4.016 8.5 66.484 ;
        RECT 3.56 4.062 8.5 66.438 ;
        RECT 3.514 4.108 8.5 66.392 ;
        RECT 3.468 4.154 8.5 66.346 ;
        RECT 3.422 4.2 8.5 66.3 ;
        RECT 3.376 4.246 8.5 66.254 ;
        RECT 3.33 4.292 8.5 66.208 ;
        RECT 3.284 4.338 8.5 66.162 ;
        RECT 3.238 4.384 8.5 66.116 ;
        RECT 3.192 4.43 8.5 66.07 ;
        RECT 3.146 4.476 8.5 66.024 ;
      LAYER MET4 ;
        RECT 0 99.5 65 107.5 ;
      LAYER MET3 ;
        RECT 0 99.5 65 107.5 ;
      LAYER MET2 ;
        RECT 0 99.5 65 107.5 ;
        RECT 45.92 78.5 57 110 ;
        RECT 8 78.5 57 89.5 ;
        RECT 33.32 78.5 44.32 110 ;
        RECT 20.66 78.5 31.66 110 ;
        RECT 8 78.5 19 110 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET5 ;
        RECT 0 68.5 65 77 ;
        RECT 0 30.788 1.5 42.212 ;
        RECT 0 30.753 1.476 42.247 ;
        RECT 0 30.707 1.43 42.293 ;
        RECT 0 30.661 1.384 42.339 ;
        RECT 0 30.615 1.338 42.385 ;
        RECT 0 30.569 1.292 42.431 ;
        RECT 0 30.523 1.246 42.477 ;
        RECT 0 30.5 1.2 42.5 ;
        RECT 0 44.288 1.5 55.712 ;
        RECT 0 44.253 1.476 55.747 ;
        RECT 0 44.207 1.43 55.793 ;
        RECT 0 44.161 1.384 55.839 ;
        RECT 0 44.115 1.338 55.885 ;
        RECT 0 44.069 1.292 55.931 ;
        RECT 0 44.023 1.246 55.977 ;
        RECT 0 44 1.2 56 ;
        RECT 0 57.788 1.5 63.212 ;
        RECT 0 57.753 1.476 63.247 ;
        RECT 0 57.707 1.43 63.293 ;
        RECT 0 57.661 1.384 63.339 ;
        RECT 0 57.615 1.338 63.385 ;
        RECT 0 57.569 1.292 63.431 ;
        RECT 0 57.523 1.246 63.477 ;
        RECT 0 57.5 1.2 63.5 ;
      LAYER MET4 ;
        RECT 0 68.5 65 77 ;
        RECT 0 30.788 1.5 42.212 ;
        RECT 0 30.753 1.476 42.247 ;
        RECT 0 30.707 1.43 42.293 ;
        RECT 0 30.661 1.384 42.339 ;
        RECT 0 30.615 1.338 42.385 ;
        RECT 0 30.569 1.292 42.431 ;
        RECT 0 30.523 1.246 42.477 ;
        RECT 0 30.5 1.2 42.5 ;
        RECT 0 44.288 1.5 55.712 ;
        RECT 0 44.253 1.476 55.747 ;
        RECT 0 44.207 1.43 55.793 ;
        RECT 0 44.161 1.384 55.839 ;
        RECT 0 44.115 1.338 55.885 ;
        RECT 0 44.069 1.292 55.931 ;
        RECT 0 44.023 1.246 55.977 ;
        RECT 0 44 1.2 56 ;
        RECT 0 57.788 1.5 63.212 ;
        RECT 0 57.753 1.476 63.247 ;
        RECT 0 57.707 1.43 63.293 ;
        RECT 0 57.661 1.384 63.339 ;
        RECT 0 57.615 1.338 63.385 ;
        RECT 0 57.569 1.292 63.431 ;
        RECT 0 57.523 1.246 63.477 ;
        RECT 0 57.5 1.2 63.5 ;
      LAYER MET3 ;
        RECT 0 68.5 65 77 ;
        RECT 0 30.788 1.5 42.212 ;
        RECT 0 30.753 1.476 42.247 ;
        RECT 0 30.707 1.43 42.293 ;
        RECT 0 30.661 1.384 42.339 ;
        RECT 0 30.615 1.338 42.385 ;
        RECT 0 30.569 1.292 42.431 ;
        RECT 0 30.523 1.246 42.477 ;
        RECT 0 30.5 1.2 42.5 ;
        RECT 0 44.288 1.5 55.712 ;
        RECT 0 44.253 1.476 55.747 ;
        RECT 0 44.207 1.43 55.793 ;
        RECT 0 44.161 1.384 55.839 ;
        RECT 0 44.115 1.338 55.885 ;
        RECT 0 44.069 1.292 55.931 ;
        RECT 0 44.023 1.246 55.977 ;
        RECT 0 44 1.2 56 ;
        RECT 0 57.788 1.5 63.212 ;
        RECT 0 57.753 1.476 63.247 ;
        RECT 0 57.707 1.43 63.293 ;
        RECT 0 57.661 1.384 63.339 ;
        RECT 0 57.615 1.338 63.385 ;
        RECT 0 57.569 1.292 63.431 ;
        RECT 0 57.523 1.246 63.477 ;
        RECT 0 57.5 1.2 63.5 ;
      LAYER MET2 ;
        RECT 0 68.5 65 77 ;
        RECT 0 57.5 65 63.5 ;
        RECT 0 44 65 56 ;
        RECT 0 30.5 65 42.5 ;
        RECT 57.015 30.5 58.205 77 ;
        RECT 51.435 30.5 52.625 77 ;
        RECT 45.855 30.5 47.045 77 ;
        RECT 40.275 30.5 41.465 77 ;
        RECT 34.695 30.5 35.885 77 ;
        RECT 29.115 30.5 30.305 77 ;
        RECT 23.535 30.5 24.725 77 ;
        RECT 17.955 30.5 19.145 77 ;
        RECT 12.375 30.5 13.565 77 ;
        RECT 6.795 30.5 7.985 77 ;
    END
  END VDDIO
  PIN VSS
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 45.25 LAYER MET2 ;
    ANTENNAPARTIALCUTAREA 6.2694 LAYER VIA4 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 1.6848 LAYER VIA2 ;
    PORT
      LAYER MET5 ;
        RECT 0 91 65 98 ;
      LAYER MET4 ;
        RECT 0 91 65 98 ;
      LAYER MET3 ;
        RECT 0 91 65 98 ;
      LAYER MET2 ;
        RECT 0 91.48 6.5 97.52 ;
        RECT 0 91.437 6.46 97.563 ;
        RECT 0 91.391 6.414 97.609 ;
        RECT 0 91.345 6.368 97.655 ;
        RECT 0 91.299 6.322 97.701 ;
        RECT 0 91.253 6.276 97.747 ;
        RECT 0 91.207 6.23 97.793 ;
        RECT 0 91.161 6.184 97.839 ;
        RECT 0 91.115 6.138 97.885 ;
        RECT 0 91.069 6.092 97.931 ;
        RECT 0 91.023 6.046 97.977 ;
        RECT 0 91 6 98 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA2 ;
    ANTENNAPARTIALCUTAREA 9.7524 LAYER VIA4 ;
    PORT
      LAYER MET5 ;
        RECT 0 78.5 65 89.5 ;
        RECT 0 3.788 1.5 15.212 ;
        RECT 0 3.753 1.476 15.247 ;
        RECT 0 3.707 1.43 15.293 ;
        RECT 0 3.661 1.384 15.339 ;
        RECT 0 3.615 1.338 15.385 ;
        RECT 0 3.569 1.292 15.431 ;
        RECT 0 3.523 1.246 15.477 ;
        RECT 0 3.5 1.2 15.5 ;
        RECT 0 17.288 1.5 28.712 ;
        RECT 0 17.253 1.476 28.747 ;
        RECT 0 17.207 1.43 28.793 ;
        RECT 0 17.161 1.384 28.839 ;
        RECT 0 17.115 1.338 28.885 ;
        RECT 0 17.069 1.292 28.931 ;
        RECT 0 17.023 1.246 28.977 ;
        RECT 0 17 1.2 29 ;
      LAYER MET4 ;
        RECT 0 78.5 65 89.5 ;
        RECT 0 3.788 1.5 15.212 ;
        RECT 0 3.753 1.476 15.247 ;
        RECT 0 3.707 1.43 15.293 ;
        RECT 0 3.661 1.384 15.339 ;
        RECT 0 3.615 1.338 15.385 ;
        RECT 0 3.569 1.292 15.431 ;
        RECT 0 3.523 1.246 15.477 ;
        RECT 0 3.5 1.2 15.5 ;
        RECT 0 17.288 1.5 28.712 ;
        RECT 0 17.253 1.476 28.747 ;
        RECT 0 17.207 1.43 28.793 ;
        RECT 0 17.161 1.384 28.839 ;
        RECT 0 17.115 1.338 28.885 ;
        RECT 0 17.069 1.292 28.931 ;
        RECT 0 17.023 1.246 28.977 ;
        RECT 0 17 1.2 29 ;
      LAYER MET3 ;
        RECT 0 78.5 65 89.5 ;
        RECT 0 3.788 1.5 15.212 ;
        RECT 0 3.753 1.476 15.247 ;
        RECT 0 3.707 1.43 15.293 ;
        RECT 0 3.661 1.384 15.339 ;
        RECT 0 3.615 1.338 15.385 ;
        RECT 0 3.569 1.292 15.431 ;
        RECT 0 3.523 1.246 15.477 ;
        RECT 0 3.5 1.2 15.5 ;
        RECT 0 17.288 1.5 28.712 ;
        RECT 0 17.253 1.476 28.747 ;
        RECT 0 17.207 1.43 28.793 ;
        RECT 0 17.161 1.384 28.839 ;
        RECT 0 17.115 1.338 28.885 ;
        RECT 0 17.069 1.292 28.931 ;
        RECT 0 17.023 1.246 28.977 ;
        RECT 0 17 1.2 29 ;
      LAYER MET2 ;
        RECT 0 17 65 29 ;
        RECT 0 3.5 65 15.5 ;
        RECT 59.805 3.5 60.995 29 ;
        RECT 54.225 3.5 55.415 29 ;
        RECT 48.645 3.5 49.835 29 ;
        RECT 43.065 3.5 44.255 29 ;
        RECT 37.485 3.5 38.675 29 ;
        RECT 31.905 3.5 33.095 29 ;
        RECT 26.325 3.5 27.515 29 ;
        RECT 20.745 3.5 21.935 29 ;
        RECT 15.165 3.5 16.355 29 ;
        RECT 9.585 3.5 10.775 29 ;
        RECT 4.005 3.5 5.195 29 ;
        RECT 0 78.98 6.5 89.02 ;
        RECT 0 78.937 6.46 89.063 ;
        RECT 0 78.891 6.414 89.109 ;
        RECT 0 78.845 6.368 89.155 ;
        RECT 0 78.799 6.322 89.201 ;
        RECT 0 78.753 6.276 89.247 ;
        RECT 0 78.707 6.23 89.293 ;
        RECT 0 78.661 6.184 89.339 ;
        RECT 0 78.615 6.138 89.385 ;
        RECT 0 78.569 6.092 89.431 ;
        RECT 0 78.523 6.046 89.477 ;
        RECT 0 78.5 6 89.5 ;
    END
  END VSSIO
  OBS
    LAYER MET1 SPACING 0.09 ;
      RECT 0 -20 65 110 ;
    LAYER MET2 SPACING 0.1 ;
      RECT 57.175 77.175 65 99.325 ;
      RECT 0 98.175 7.825 99.325 ;
      RECT 6.675 77.175 7.825 99.325 ;
      RECT 6.175 98.152 7.825 99.325 ;
      RECT 6.635 97.695 7.825 99.325 ;
      RECT 6.221 98.106 7.825 99.325 ;
      RECT 6.589 97.738 7.825 99.325 ;
      RECT 6.267 98.06 7.825 99.325 ;
      RECT 6.543 97.784 7.825 99.325 ;
      RECT 6.313 98.014 7.825 99.325 ;
      RECT 6.497 97.83 7.825 99.325 ;
      RECT 6.359 97.968 7.825 99.325 ;
      RECT 6.451 97.876 7.825 99.325 ;
      RECT 6.405 97.922 7.825 99.325 ;
      RECT 6.635 89.195 7.825 91.305 ;
      RECT 6.589 89.238 7.825 91.262 ;
      RECT 6.543 89.284 7.825 91.216 ;
      RECT 6.497 89.33 7.825 91.17 ;
      RECT 6.451 89.376 7.825 91.124 ;
      RECT 6.405 89.422 7.825 91.078 ;
      RECT 6.359 89.468 7.825 91.032 ;
      RECT 6.313 89.514 7.825 90.986 ;
      RECT 6.267 89.56 7.825 90.94 ;
      RECT 6.221 89.606 7.825 90.894 ;
      RECT 6.175 89.652 7.825 90.848 ;
      RECT 0 89.675 7.825 90.825 ;
      RECT 6.635 77.175 7.825 78.805 ;
      RECT 6.589 77.175 7.825 78.762 ;
      RECT 6.543 77.175 7.825 78.716 ;
      RECT 6.497 77.175 7.825 78.67 ;
      RECT 6.451 77.175 7.825 78.624 ;
      RECT 6.405 77.175 7.825 78.578 ;
      RECT 6.359 77.175 7.825 78.532 ;
      RECT 6.313 77.175 7.825 78.486 ;
      RECT 6.267 77.175 7.825 78.44 ;
      RECT 6.221 77.175 7.825 78.394 ;
      RECT 6.175 77.175 7.825 78.348 ;
      RECT 0 77.175 65 78.325 ;
      RECT 0 -20 65 3.325 ;
      RECT 61.17 15.675 65 16.825 ;
      RECT 0 29.175 65 30.325 ;
      RECT 58.38 42.675 65 43.825 ;
      RECT 58.38 56.175 65 57.325 ;
      RECT 58.38 63.675 65 68.325 ;
      RECT 57.175 107.675 65 110 ;
      RECT 55.59 15.675 59.63 16.825 ;
      RECT 52.8 42.675 56.84 43.825 ;
      RECT 52.8 56.175 56.84 57.325 ;
      RECT 52.8 63.675 56.84 68.325 ;
      RECT 50.01 15.675 54.05 16.825 ;
      RECT 47.22 42.675 51.26 43.825 ;
      RECT 47.22 56.175 51.26 57.325 ;
      RECT 47.22 63.675 51.26 68.325 ;
      RECT 44.43 15.675 48.47 16.825 ;
      RECT 44.495 89.675 45.745 99.325 ;
      RECT 41.64 42.675 45.68 43.825 ;
      RECT 41.64 56.175 45.68 57.325 ;
      RECT 41.64 63.675 45.68 68.325 ;
      RECT 38.85 15.675 42.89 16.825 ;
      RECT 36.06 42.675 40.1 43.825 ;
      RECT 36.06 56.175 40.1 57.325 ;
      RECT 36.06 63.675 40.1 68.325 ;
      RECT 33.27 15.675 37.31 16.825 ;
      RECT 30.48 42.675 34.52 43.825 ;
      RECT 30.48 56.175 34.52 57.325 ;
      RECT 30.48 63.675 34.52 68.325 ;
      RECT 31.835 89.675 33.145 99.325 ;
      RECT 27.69 15.675 31.73 16.825 ;
      RECT 24.9 42.675 28.94 43.825 ;
      RECT 24.9 56.175 28.94 57.325 ;
      RECT 24.9 63.675 28.94 68.325 ;
      RECT 22.11 15.675 26.15 16.825 ;
      RECT 19.32 42.675 23.36 43.825 ;
      RECT 19.32 56.175 23.36 57.325 ;
      RECT 19.32 63.675 23.36 68.325 ;
      RECT 16.53 15.675 20.57 16.825 ;
      RECT 19.175 89.675 20.485 99.325 ;
      RECT 13.74 42.675 17.78 43.825 ;
      RECT 13.74 56.175 17.78 57.325 ;
      RECT 13.74 63.675 17.78 68.325 ;
      RECT 10.95 15.675 14.99 16.825 ;
      RECT 8.16 42.675 12.2 43.825 ;
      RECT 8.16 56.175 12.2 57.325 ;
      RECT 8.16 63.675 12.2 68.325 ;
      RECT 5.37 15.675 9.41 16.825 ;
      RECT 0 107.675 7.825 110 ;
      RECT 0 42.675 6.62 43.825 ;
      RECT 0 56.175 6.62 57.325 ;
      RECT 0 63.675 6.62 68.325 ;
      RECT 0 15.675 3.83 16.825 ;
    LAYER MET3 SPACING 0.1 ;
      RECT 62 63.665 65 68.325 ;
      RECT 58.37 -20 61 68.325 ;
      RECT 52.79 57.5 56.85 68.325 ;
      RECT 47.21 57.5 51.27 68.325 ;
      RECT 41.63 57.5 45.69 68.325 ;
      RECT 36.05 57.5 40.11 68.325 ;
      RECT 30.47 -20 34.53 68.325 ;
      RECT 24.89 57.5 28.95 68.325 ;
      RECT 19.31 57.5 23.37 68.325 ;
      RECT 13.73 57.5 17.79 68.325 ;
      RECT 8.15 57.5 12.21 68.325 ;
      RECT 4 -20 6.63 68.325 ;
      RECT 0 63.675 3 68.325 ;
      RECT 1.375 63.665 3 68.325 ;
      RECT 4 57.5 61 67 ;
      RECT 57 -20 61 67 ;
      RECT 43 -20 50.5 67 ;
      RECT 29 -20 36.5 67 ;
      RECT 15 -20 22.5 67 ;
      RECT 4 -20 8.5 67 ;
      RECT 62 56.165 65 57.335 ;
      RECT 41.63 56.165 51.27 57.335 ;
      RECT 24.89 56.165 40.11 57.335 ;
      RECT 13.73 56.165 23.37 57.335 ;
      RECT 4 56.165 12.21 57.335 ;
      RECT 1.375 56.165 3 57.335 ;
      RECT 0 56.175 3 57.325 ;
      RECT 4 43.5 61 51 ;
      RECT 62 42.665 65 43.835 ;
      RECT 1.375 42.665 3 43.835 ;
      RECT 0 42.675 3 43.825 ;
      RECT 52.79 42.665 56.85 51 ;
      RECT 41.63 42.665 51.27 51 ;
      RECT 24.89 42.665 40.11 51 ;
      RECT 13.73 42.665 23.37 51 ;
      RECT 4 42.665 12.21 51 ;
      RECT 4 29.165 61 37 ;
      RECT 62 29.165 65 30.335 ;
      RECT 1.375 29.165 3 30.335 ;
      RECT 0 29.175 3 30.325 ;
      RECT 4 15.5 61 23 ;
      RECT 62 15.665 65 16.835 ;
      RECT 1.375 15.665 3 16.835 ;
      RECT 0 15.675 3 16.825 ;
      RECT 4 -20 61 9 ;
      RECT 1.375 -20 65 3.335 ;
      RECT 0 -20 65 3.325 ;
      RECT 61.966 4.483 62 68.325 ;
      RECT 61.92 4.443 61.966 68.325 ;
      RECT 61.874 4.397 61.92 68.325 ;
      RECT 61.828 4.351 61.874 68.325 ;
      RECT 61.782 4.305 61.828 68.325 ;
      RECT 61.736 4.259 61.782 68.325 ;
      RECT 61.69 4.213 61.736 68.325 ;
      RECT 61.644 4.167 61.69 68.325 ;
      RECT 61.598 4.121 61.644 68.325 ;
      RECT 61.552 4.075 61.598 68.325 ;
      RECT 61.506 4.029 61.552 68.325 ;
      RECT 61.46 3.983 61.506 68.325 ;
      RECT 61.414 3.937 61.46 68.325 ;
      RECT 61.368 3.891 61.414 68.325 ;
      RECT 61.322 3.845 61.368 68.325 ;
      RECT 61.276 3.799 61.322 68.325 ;
      RECT 61.23 3.753 61.276 68.325 ;
      RECT 61.184 3.707 61.23 68.325 ;
      RECT 61.138 3.661 61.184 68.325 ;
      RECT 61.092 3.615 61.138 68.325 ;
      RECT 61.046 3.569 61.092 68.325 ;
      RECT 61 3.523 61.046 68.325 ;
      RECT 3.966 3.517 4 68.325 ;
      RECT 3.92 3.557 3.966 68.325 ;
      RECT 3.874 3.603 3.92 68.325 ;
      RECT 3.828 3.649 3.874 68.325 ;
      RECT 3.782 3.695 3.828 68.325 ;
      RECT 3.736 3.741 3.782 68.325 ;
      RECT 3.69 3.787 3.736 68.325 ;
      RECT 3.644 3.833 3.69 68.325 ;
      RECT 3.598 3.879 3.644 68.325 ;
      RECT 3.552 3.925 3.598 68.325 ;
      RECT 3.506 3.971 3.552 68.325 ;
      RECT 3.46 4.017 3.506 68.325 ;
      RECT 3.414 4.063 3.46 68.325 ;
      RECT 3.368 4.109 3.414 68.325 ;
      RECT 3.322 4.155 3.368 68.325 ;
      RECT 3.276 4.201 3.322 68.325 ;
      RECT 3.23 4.247 3.276 68.325 ;
      RECT 3.184 4.293 3.23 68.325 ;
      RECT 3.138 4.339 3.184 68.325 ;
      RECT 3.092 4.385 3.138 68.325 ;
      RECT 3.046 4.431 3.092 68.325 ;
      RECT 3 4.477 3.046 68.325 ;
      RECT 63.8 3.5 65 15.5 ;
      RECT 63.776 3.512 65 15.488 ;
      RECT 63.73 3.547 65 15.453 ;
      RECT 63.684 3.593 65 15.407 ;
      RECT 63.638 3.639 65 15.361 ;
      RECT 63.592 3.685 65 15.315 ;
      RECT 63.546 3.731 65 15.269 ;
      RECT 63.5 3.777 65 15.223 ;
      RECT 63.8 17 65 29 ;
      RECT 63.776 17.012 65 28.988 ;
      RECT 63.73 17.047 65 28.953 ;
      RECT 63.684 17.093 65 28.907 ;
      RECT 63.638 17.139 65 28.861 ;
      RECT 63.592 17.185 65 28.815 ;
      RECT 63.546 17.231 65 28.769 ;
      RECT 63.5 17.277 65 28.723 ;
      RECT 63.8 30.5 65 42.5 ;
      RECT 63.776 30.512 65 42.488 ;
      RECT 63.73 30.547 65 42.453 ;
      RECT 63.684 30.593 65 42.407 ;
      RECT 63.638 30.639 65 42.361 ;
      RECT 63.592 30.685 65 42.315 ;
      RECT 63.546 30.731 65 42.269 ;
      RECT 63.5 30.777 65 42.223 ;
      RECT 63.8 44 65 56 ;
      RECT 63.776 44.012 65 55.988 ;
      RECT 63.73 44.047 65 55.953 ;
      RECT 63.684 44.093 65 55.907 ;
      RECT 63.638 44.139 65 55.861 ;
      RECT 63.592 44.185 65 55.815 ;
      RECT 63.546 44.231 65 55.769 ;
      RECT 63.5 44.277 65 55.723 ;
      RECT 63.8 57.5 65 63.5 ;
      RECT 63.776 57.512 65 63.488 ;
      RECT 63.73 57.547 65 63.453 ;
      RECT 63.684 57.593 65 63.407 ;
      RECT 63.638 57.639 65 63.361 ;
      RECT 63.592 57.685 65 63.315 ;
      RECT 63.546 57.731 65 63.269 ;
      RECT 63.5 57.777 65 63.223 ;
      RECT 57.175 107.675 65 110 ;
      RECT 57.165 107.675 65 108.825 ;
      RECT 0 107.675 7.825 110 ;
      RECT 0 107.675 7.835 108.825 ;
      RECT 0 77.175 65 78.325 ;
      RECT 57.165 89.675 65 90.825 ;
      RECT 57.165 98.175 65 99.325 ;
      RECT 52.79 56.165 56.85 57.335 ;
      RECT 44.485 89.675 45.755 90.825 ;
      RECT 44.485 98.175 45.755 99.325 ;
      RECT 31.825 89.675 33.155 90.825 ;
      RECT 31.825 98.175 33.155 99.325 ;
      RECT 19.165 89.675 20.495 90.825 ;
      RECT 19.165 98.175 20.495 99.325 ;
      RECT 0 89.675 7.835 90.825 ;
      RECT 0 98.175 7.835 99.325 ;
    LAYER MET4 SPACING 0.1 ;
      RECT 0 63.675 65 68.325 ;
      RECT 1.675 -20 65 68.325 ;
      RECT 1.375 63.652 65 68.325 ;
      RECT 1.651 63.387 65 68.325 ;
      RECT 1.421 63.606 65 68.325 ;
      RECT 1.605 63.422 65 68.325 ;
      RECT 1.467 63.56 65 68.325 ;
      RECT 1.559 63.468 65 68.325 ;
      RECT 1.513 63.514 65 68.325 ;
      RECT 1.651 55.887 65 57.613 ;
      RECT 1.605 55.922 65 57.578 ;
      RECT 1.559 55.968 65 57.532 ;
      RECT 1.513 56.014 65 57.486 ;
      RECT 1.467 56.06 65 57.44 ;
      RECT 1.421 56.106 65 57.394 ;
      RECT 1.375 56.152 65 57.348 ;
      RECT 0 56.175 65 57.325 ;
      RECT 1.651 42.387 65 44.113 ;
      RECT 1.605 42.422 65 44.078 ;
      RECT 1.559 42.468 65 44.032 ;
      RECT 1.513 42.514 65 43.986 ;
      RECT 1.467 42.56 65 43.94 ;
      RECT 1.421 42.606 65 43.894 ;
      RECT 1.375 42.652 65 43.848 ;
      RECT 0 42.675 65 43.825 ;
      RECT 1.651 28.887 65 30.613 ;
      RECT 1.605 28.922 65 30.578 ;
      RECT 1.559 28.968 65 30.532 ;
      RECT 1.513 29.014 65 30.486 ;
      RECT 1.467 29.06 65 30.44 ;
      RECT 1.421 29.106 65 30.394 ;
      RECT 1.375 29.152 65 30.348 ;
      RECT 0 29.175 65 30.325 ;
      RECT 1.651 15.387 65 17.113 ;
      RECT 1.605 15.422 65 17.078 ;
      RECT 1.559 15.468 65 17.032 ;
      RECT 1.513 15.514 65 16.986 ;
      RECT 1.467 15.56 65 16.94 ;
      RECT 1.421 15.606 65 16.894 ;
      RECT 1.375 15.652 65 16.848 ;
      RECT 0 15.675 65 16.825 ;
      RECT 1.651 -20 65 3.613 ;
      RECT 1.605 -20 65 3.578 ;
      RECT 1.559 -20 65 3.532 ;
      RECT 1.513 -20 65 3.486 ;
      RECT 1.467 -20 65 3.44 ;
      RECT 1.421 -20 65 3.394 ;
      RECT 1.375 -20 65 3.348 ;
      RECT 0 -20 65 3.325 ;
      RECT 57.175 107.675 65 110 ;
      RECT 0 107.675 7.825 110 ;
      RECT 0 107.675 65 108.825 ;
      RECT 0 77.175 65 78.325 ;
      RECT 0 89.675 65 90.825 ;
      RECT 0 98.175 65 99.325 ;
    LAYER MET5 SPACING 0.1 ;
      RECT 0 63.83 65 68.17 ;
      RECT 1.83 -20 65 68.17 ;
      RECT 1.53 63.807 65 68.17 ;
      RECT 1.806 63.542 65 68.17 ;
      RECT 1.576 63.761 65 68.17 ;
      RECT 1.76 63.577 65 68.17 ;
      RECT 1.622 63.715 65 68.17 ;
      RECT 1.714 63.623 65 68.17 ;
      RECT 1.668 63.669 65 68.17 ;
      RECT 1.806 56.042 65 57.458 ;
      RECT 1.76 56.077 65 57.423 ;
      RECT 1.714 56.123 65 57.377 ;
      RECT 1.668 56.169 65 57.331 ;
      RECT 1.622 56.215 65 57.285 ;
      RECT 1.576 56.261 65 57.239 ;
      RECT 1.53 56.307 65 57.193 ;
      RECT 0 56.33 65 57.17 ;
      RECT 1.806 42.542 65 43.958 ;
      RECT 1.76 42.577 65 43.923 ;
      RECT 1.714 42.623 65 43.877 ;
      RECT 1.668 42.669 65 43.831 ;
      RECT 1.622 42.715 65 43.785 ;
      RECT 1.576 42.761 65 43.739 ;
      RECT 1.53 42.807 65 43.693 ;
      RECT 0 42.83 65 43.67 ;
      RECT 1.806 29.042 65 30.458 ;
      RECT 1.76 29.077 65 30.423 ;
      RECT 1.714 29.123 65 30.377 ;
      RECT 1.668 29.169 65 30.331 ;
      RECT 1.622 29.215 65 30.285 ;
      RECT 1.576 29.261 65 30.239 ;
      RECT 1.53 29.307 65 30.193 ;
      RECT 0 29.33 65 30.17 ;
      RECT 1.806 15.542 65 16.958 ;
      RECT 1.76 15.577 65 16.923 ;
      RECT 1.714 15.623 65 16.877 ;
      RECT 1.668 15.669 65 16.831 ;
      RECT 1.622 15.715 65 16.785 ;
      RECT 1.576 15.761 65 16.739 ;
      RECT 1.53 15.807 65 16.693 ;
      RECT 0 15.83 65 16.67 ;
      RECT 1.806 -20 65 3.458 ;
      RECT 1.76 -20 65 3.423 ;
      RECT 1.714 -20 65 3.377 ;
      RECT 1.668 -20 65 3.331 ;
      RECT 1.622 -20 65 3.285 ;
      RECT 1.576 -20 65 3.239 ;
      RECT 1.53 -20 65 3.193 ;
      RECT 0 -20 65 3.17 ;
      RECT 57.33 107.83 65 110 ;
      RECT 0 107.83 7.67 110 ;
      RECT 0 107.83 65 108.67 ;
      RECT 0 77.33 65 78.17 ;
      RECT 0 89.83 65 90.67 ;
      RECT 0 98.33 65 99.17 ;
    LAYER T4M2 SPACING 0.4 ;
      RECT 64.585 -20 65 0.453 ;
      RECT 0 -20 0.436 0.432 ;
      RECT 64.539 -20 65 0.407 ;
      RECT 0 -20 0.482 0.386 ;
      RECT 64.493 -20 65 0.361 ;
      RECT 0 -20 0.528 0.34 ;
      RECT 64.447 -20 65 0.315 ;
      RECT 0 -20 0.574 0.294 ;
      RECT 64.401 -20 65 0.269 ;
      RECT 0 -20 0.62 0.248 ;
      RECT 64.355 -20 65 0.223 ;
      RECT 0 -20 0.645 0.212 ;
      RECT 64.346 -20 65 0.195 ;
      RECT 0 -20 0.691 0.177 ;
      RECT 64.3 -20 65 0.168 ;
      RECT 0 -20 0.7 0.149 ;
      RECT 0 -20 65 -3.3 ;
      RECT 57.6 108.1 65 110 ;
      RECT 0 108.1 7.4 110 ;
    LAYER RDL SPACING 2 ;
      RECT 0 -20 65 -4.9 ;
      RECT 0 71.9 65 110 ;
      RECT 3 4.5 62 63.5 ;
  END
END P65_1233_VDD3

MACRO P65_1233_VDDIO3
  CLASS PAD ;
  ORIGIN 0 20 ;
  FOREIGN P65_1233_VDDIO3 0 -20 ;
  SIZE 65 BY 130 ;
  SYMMETRY X Y R90 ;
  SITE IOSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET4 ;
        RECT 0 100.483 6.5 106.517 ;
        RECT 0 100.443 6.466 106.557 ;
        RECT 0 100.397 6.42 106.603 ;
        RECT 0 100.351 6.374 106.649 ;
        RECT 0 100.305 6.328 106.695 ;
        RECT 0 100.259 6.282 106.741 ;
        RECT 0 100.213 6.236 106.787 ;
        RECT 0 100.167 6.19 106.833 ;
        RECT 0 100.121 6.144 106.879 ;
        RECT 0 100.075 6.098 106.925 ;
        RECT 0 100.029 6.052 106.971 ;
        RECT 0 99.983 6.006 107.017 ;
        RECT 0 99.937 5.96 107.063 ;
        RECT 0 99.891 5.914 107.109 ;
        RECT 0 99.845 5.868 107.155 ;
        RECT 0 99.799 5.822 107.201 ;
        RECT 0 99.753 5.776 107.247 ;
        RECT 0 99.707 5.73 107.293 ;
        RECT 0 99.661 5.684 107.339 ;
        RECT 0 99.615 5.638 107.385 ;
        RECT 0 99.569 5.592 107.431 ;
        RECT 0 99.523 5.546 107.477 ;
        RECT 0 99.5 5.5 107.5 ;
      LAYER MET3 ;
        RECT 0 100.483 6.5 106.517 ;
        RECT 0 100.443 6.466 106.557 ;
        RECT 0 100.397 6.42 106.603 ;
        RECT 0 100.351 6.374 106.649 ;
        RECT 0 100.305 6.328 106.695 ;
        RECT 0 100.259 6.282 106.741 ;
        RECT 0 100.213 6.236 106.787 ;
        RECT 0 100.167 6.19 106.833 ;
        RECT 0 100.121 6.144 106.879 ;
        RECT 0 100.075 6.098 106.925 ;
        RECT 0 100.029 6.052 106.971 ;
        RECT 0 99.983 6.006 107.017 ;
        RECT 0 99.937 5.96 107.063 ;
        RECT 0 99.891 5.914 107.109 ;
        RECT 0 99.845 5.868 107.155 ;
        RECT 0 99.799 5.822 107.201 ;
        RECT 0 99.753 5.776 107.247 ;
        RECT 0 99.707 5.73 107.293 ;
        RECT 0 99.661 5.684 107.339 ;
        RECT 0 99.615 5.638 107.385 ;
        RECT 0 99.569 5.592 107.431 ;
        RECT 0 99.523 5.546 107.477 ;
        RECT 0 99.5 5.5 107.5 ;
    END
    PORT
      CLASS CORE ;
      LAYER MET5 ;
        RECT 0 99.5 65 107.5 ;
      LAYER MET2 ;
        RECT 0 99.5 65 107.5 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET5 ;
        RECT 0 68.5 65 77 ;
        RECT 57 57.5 65 63.5 ;
        RECT 57 44 65 56 ;
        RECT 57 30.5 65 42.5 ;
        RECT 57 4.483 62 63.5 ;
        RECT 57 4.443 61.966 63.5 ;
        RECT 3.046 4.431 61.92 12 ;
        RECT 57 4.397 61.92 63.5 ;
        RECT 3.092 4.385 61.874 12 ;
        RECT 57 4.351 61.874 63.5 ;
        RECT 3.138 4.339 61.828 12 ;
        RECT 57 4.305 61.828 63.5 ;
        RECT 3.184 4.293 61.782 12 ;
        RECT 57 4.259 61.782 63.5 ;
        RECT 3.23 4.247 61.736 12 ;
        RECT 57 4.213 61.736 63.5 ;
        RECT 3.276 4.201 61.69 12 ;
        RECT 57 4.167 61.69 63.5 ;
        RECT 3.322 4.155 61.644 12 ;
        RECT 57 4.121 61.644 63.5 ;
        RECT 3.368 4.109 61.598 12 ;
        RECT 57 4.075 61.598 63.5 ;
        RECT 3.414 4.063 61.552 12 ;
        RECT 57 4.029 61.552 63.5 ;
        RECT 3.46 4.017 61.506 12 ;
        RECT 57 3.983 61.506 63.5 ;
        RECT 3.506 3.971 61.46 12 ;
        RECT 57 3.937 61.46 63.5 ;
        RECT 3.552 3.925 61.414 12 ;
        RECT 57 3.891 61.414 63.5 ;
        RECT 3.598 3.879 61.368 12 ;
        RECT 57 3.845 61.368 63.5 ;
        RECT 3.644 3.833 61.322 12 ;
        RECT 57 3.799 61.322 63.5 ;
        RECT 3.69 3.787 61.276 12 ;
        RECT 57 3.753 61.276 63.5 ;
        RECT 3.736 3.741 61.23 12 ;
        RECT 57 3.707 61.23 63.5 ;
        RECT 3.782 3.695 61.184 12 ;
        RECT 57 3.661 61.184 63.5 ;
        RECT 3.828 3.649 61.138 12 ;
        RECT 57 3.615 61.138 63.5 ;
        RECT 3.874 3.603 61.092 12 ;
        RECT 57 3.569 61.092 63.5 ;
        RECT 3.92 3.557 61.046 12 ;
        RECT 57 3.523 61.046 63.5 ;
        RECT 3.966 3.517 61 12 ;
        RECT 46 61.08 58 77 ;
        RECT 0 47.08 65 54.58 ;
        RECT 0 33.08 65 40.58 ;
        RECT 3 19.08 62 26.58 ;
        RECT 4 0 61 12 ;
        RECT 43 0 50.5 63.5 ;
        RECT 33.27 61.08 44.34 77 ;
        RECT 29 0 36.5 63.5 ;
        RECT 20.66 61.08 31.66 77 ;
        RECT 15 0 22.5 63.5 ;
        RECT 7 61.08 19 77 ;
        RECT 0 57.5 8.5 63.5 ;
        RECT 3 4.477 8.5 63.5 ;
        RECT 0 44 8.5 56 ;
        RECT 0 30.5 8.5 42.5 ;
        RECT 8 109 57 110 ;
      LAYER T4M2 ;
        RECT 3.1 57.4 61.9 76.9 ;
        RECT 57 4.528 61.9 76.9 ;
        RECT 57 4.488 61.866 76.9 ;
        RECT 3.146 4.471 61.82 8.9 ;
        RECT 57 4.442 61.82 76.9 ;
        RECT 3.192 4.425 61.774 8.9 ;
        RECT 57 4.396 61.774 76.9 ;
        RECT 3.238 4.379 61.728 8.9 ;
        RECT 57 4.35 61.728 76.9 ;
        RECT 3.284 4.333 61.682 8.9 ;
        RECT 57 4.304 61.682 76.9 ;
        RECT 3.33 4.287 61.636 8.9 ;
        RECT 57 4.258 61.636 76.9 ;
        RECT 3.376 4.241 61.59 8.9 ;
        RECT 57 4.212 61.59 76.9 ;
        RECT 3.422 4.195 61.544 8.9 ;
        RECT 57 4.166 61.544 76.9 ;
        RECT 3.468 4.149 61.498 8.9 ;
        RECT 57 4.12 61.498 76.9 ;
        RECT 3.514 4.103 61.452 8.9 ;
        RECT 57 4.074 61.452 76.9 ;
        RECT 3.56 4.057 61.406 8.9 ;
        RECT 57 4.028 61.406 76.9 ;
        RECT 3.606 4.011 61.36 8.9 ;
        RECT 57 3.982 61.36 76.9 ;
        RECT 3.652 3.965 61.314 8.9 ;
        RECT 57 3.936 61.314 76.9 ;
        RECT 3.698 3.919 61.268 8.9 ;
        RECT 57 3.89 61.268 76.9 ;
        RECT 3.744 3.873 61.222 8.9 ;
        RECT 57 3.844 61.222 76.9 ;
        RECT 3.79 3.827 61.176 8.9 ;
        RECT 57 3.798 61.176 76.9 ;
        RECT 3.836 3.781 61.13 8.9 ;
        RECT 57 3.752 61.13 76.9 ;
        RECT 3.882 3.735 61.084 8.9 ;
        RECT 57 3.706 61.084 76.9 ;
        RECT 3.928 3.689 61.038 8.9 ;
        RECT 57 3.66 61.038 76.9 ;
        RECT 3.974 3.643 60.992 8.9 ;
        RECT 57 3.614 60.992 76.9 ;
        RECT 4.02 3.597 60.946 8.9 ;
        RECT 57 3.568 60.946 76.9 ;
        RECT 4.066 3.557 60.9 8.9 ;
        RECT 3.1 43.4 61.9 50.9 ;
        RECT 3.1 29.4 61.9 36.9 ;
        RECT 3.1 15.4 61.9 22.9 ;
        RECT 4.1 0.1 60.9 8.9 ;
        RECT 43 0.1 50.5 76.9 ;
        RECT 29 0.1 36.5 76.9 ;
        RECT 15 0.1 22.5 76.9 ;
        RECT 3.1 4.517 8.5 76.9 ;
      LAYER MET4 ;
        RECT 0 68.5 65 77 ;
        RECT 57 57.5 65 63.5 ;
        RECT 57 44 65 56 ;
        RECT 57 30.5 65 42.5 ;
        RECT 57 4.483 62 63.5 ;
        RECT 57 4.443 61.966 63.5 ;
        RECT 3.046 4.431 61.92 12 ;
        RECT 57 4.397 61.92 63.5 ;
        RECT 3.092 4.385 61.874 12 ;
        RECT 57 4.351 61.874 63.5 ;
        RECT 3.138 4.339 61.828 12 ;
        RECT 57 4.305 61.828 63.5 ;
        RECT 3.184 4.293 61.782 12 ;
        RECT 57 4.259 61.782 63.5 ;
        RECT 3.23 4.247 61.736 12 ;
        RECT 57 4.213 61.736 63.5 ;
        RECT 3.276 4.201 61.69 12 ;
        RECT 57 4.167 61.69 63.5 ;
        RECT 3.322 4.155 61.644 12 ;
        RECT 57 4.121 61.644 63.5 ;
        RECT 3.368 4.109 61.598 12 ;
        RECT 57 4.075 61.598 63.5 ;
        RECT 3.414 4.063 61.552 12 ;
        RECT 57 4.029 61.552 63.5 ;
        RECT 3.46 4.017 61.506 12 ;
        RECT 57 3.983 61.506 63.5 ;
        RECT 3.506 3.971 61.46 12 ;
        RECT 57 3.937 61.46 63.5 ;
        RECT 3.552 3.925 61.414 12 ;
        RECT 57 3.891 61.414 63.5 ;
        RECT 3.598 3.879 61.368 12 ;
        RECT 57 3.845 61.368 63.5 ;
        RECT 3.644 3.833 61.322 12 ;
        RECT 57 3.799 61.322 63.5 ;
        RECT 3.69 3.787 61.276 12 ;
        RECT 57 3.753 61.276 63.5 ;
        RECT 3.736 3.741 61.23 12 ;
        RECT 57 3.707 61.23 63.5 ;
        RECT 3.782 3.695 61.184 12 ;
        RECT 57 3.661 61.184 63.5 ;
        RECT 3.828 3.649 61.138 12 ;
        RECT 57 3.615 61.138 63.5 ;
        RECT 3.874 3.603 61.092 12 ;
        RECT 57 3.569 61.092 63.5 ;
        RECT 3.92 3.557 61.046 12 ;
        RECT 57 3.523 61.046 63.5 ;
        RECT 3.966 3.517 61 12 ;
        RECT 46 61.08 58 77 ;
        RECT 8 109 57 110 ;
        RECT 46 61.08 57 110 ;
        RECT 0 47.08 65 54.58 ;
        RECT 0 33.08 65 40.58 ;
        RECT 3 19.08 62 26.58 ;
        RECT 4 0 61 12 ;
        RECT 43 0 50.5 63.5 ;
        RECT 33.27 61.08 44.34 110 ;
        RECT 29 0 36.5 63.5 ;
        RECT 20.66 61.08 31.66 110 ;
        RECT 15 0 22.5 63.5 ;
        RECT 8 61.08 19 110 ;
        RECT 0 57.5 8.5 63.5 ;
        RECT 7 61.08 19 77 ;
        RECT 3 4.477 8.5 63.5 ;
        RECT 0 44 8.5 56 ;
        RECT 0 30.5 8.5 42.5 ;
      LAYER MET3 ;
        RECT 0 68.5 65 77 ;
        RECT 57 57.5 65 63.5 ;
        RECT 57 44 65 56 ;
        RECT 57 30.5 65 42.5 ;
        RECT 57 4.483 62 63.5 ;
        RECT 57 4.443 61.966 63.5 ;
        RECT 3.046 4.431 61.92 12 ;
        RECT 57 4.397 61.92 63.5 ;
        RECT 3.092 4.385 61.874 12 ;
        RECT 57 4.351 61.874 63.5 ;
        RECT 3.138 4.339 61.828 12 ;
        RECT 57 4.305 61.828 63.5 ;
        RECT 3.184 4.293 61.782 12 ;
        RECT 57 4.259 61.782 63.5 ;
        RECT 3.23 4.247 61.736 12 ;
        RECT 57 4.213 61.736 63.5 ;
        RECT 3.276 4.201 61.69 12 ;
        RECT 57 4.167 61.69 63.5 ;
        RECT 3.322 4.155 61.644 12 ;
        RECT 57 4.121 61.644 63.5 ;
        RECT 3.368 4.109 61.598 12 ;
        RECT 57 4.075 61.598 63.5 ;
        RECT 3.414 4.063 61.552 12 ;
        RECT 57 4.029 61.552 63.5 ;
        RECT 3.46 4.017 61.506 12 ;
        RECT 57 3.983 61.506 63.5 ;
        RECT 3.506 3.971 61.46 12 ;
        RECT 57 3.937 61.46 63.5 ;
        RECT 3.552 3.925 61.414 12 ;
        RECT 57 3.891 61.414 63.5 ;
        RECT 3.598 3.879 61.368 12 ;
        RECT 57 3.845 61.368 63.5 ;
        RECT 3.644 3.833 61.322 12 ;
        RECT 57 3.799 61.322 63.5 ;
        RECT 3.69 3.787 61.276 12 ;
        RECT 57 3.753 61.276 63.5 ;
        RECT 3.736 3.741 61.23 12 ;
        RECT 57 3.707 61.23 63.5 ;
        RECT 3.782 3.695 61.184 12 ;
        RECT 57 3.661 61.184 63.5 ;
        RECT 3.828 3.649 61.138 12 ;
        RECT 57 3.615 61.138 63.5 ;
        RECT 3.874 3.603 61.092 12 ;
        RECT 57 3.569 61.092 63.5 ;
        RECT 3.92 3.557 61.046 12 ;
        RECT 57 3.523 61.046 63.5 ;
        RECT 3.966 3.517 61 12 ;
        RECT 46 61.08 58 77 ;
        RECT 8 109 57 110 ;
        RECT 46 61.08 57 110 ;
        RECT 0 47.08 65 54.58 ;
        RECT 0 33.08 65 40.58 ;
        RECT 3 19.08 62 26.58 ;
        RECT 4 0 61 12 ;
        RECT 43 0 50.5 63.5 ;
        RECT 33.27 61.08 44.34 110 ;
        RECT 29 0 36.5 63.5 ;
        RECT 20.66 61.08 31.66 110 ;
        RECT 15 0 22.5 63.5 ;
        RECT 8 61.08 19 110 ;
        RECT 0 57.5 8.5 63.5 ;
        RECT 7 61.08 19 77 ;
        RECT 3 4.477 8.5 63.5 ;
        RECT 0 44 8.5 56 ;
        RECT 0 30.5 8.5 42.5 ;
      LAYER MET2 ;
        RECT 0 57.5 65 63.5 ;
        RECT 0 44 65 56 ;
        RECT 0 30.5 65 42.5 ;
        RECT 56.015 30.5 59.205 63.5 ;
        RECT 50.435 30.5 53.625 63.5 ;
        RECT 44.855 30.5 48.045 63.5 ;
        RECT 39.275 30.5 42.465 63.5 ;
        RECT 33.695 30.5 36.885 63.5 ;
        RECT 28.115 30.5 31.305 63.5 ;
        RECT 22.535 30.5 25.725 63.5 ;
        RECT 16.955 30.5 20.145 63.5 ;
        RECT 11.375 30.5 14.565 63.5 ;
        RECT 5.795 30.5 8.985 63.5 ;
        RECT 0 68.5 65 77 ;
        RECT 8 109 57 110 ;
    END
  END VDDIO
  PIN VSS
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 44.5 LAYER MET4 ;
    ANTENNAPARTIALMETALAREA 44.5 LAYER MET3 ;
    ANTENNAPARTIALCUTAREA 1.053 LAYER VIA4 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 4.617 LAYER VIA2 ;
    PORT
      LAYER MET5 ;
        RECT 0 91 65 98 ;
      LAYER MET4 ;
        RECT 0 91.983 6.5 97.017 ;
        RECT 0 91.943 6.466 97.057 ;
        RECT 0 91.897 6.42 97.103 ;
        RECT 0 91.851 6.374 97.149 ;
        RECT 0 91.805 6.328 97.195 ;
        RECT 0 91.759 6.282 97.241 ;
        RECT 0 91.713 6.236 97.287 ;
        RECT 0 91.667 6.19 97.333 ;
        RECT 0 91.621 6.144 97.379 ;
        RECT 0 91.575 6.098 97.425 ;
        RECT 0 91.529 6.052 97.471 ;
        RECT 0 91.483 6.006 97.517 ;
        RECT 0 91.437 5.96 97.563 ;
        RECT 0 91.391 5.914 97.609 ;
        RECT 0 91.345 5.868 97.655 ;
        RECT 0 91.299 5.822 97.701 ;
        RECT 0 91.253 5.776 97.747 ;
        RECT 0 91.207 5.73 97.793 ;
        RECT 0 91.161 5.684 97.839 ;
        RECT 0 91.115 5.638 97.885 ;
        RECT 0 91.069 5.592 97.931 ;
        RECT 0 91.023 5.546 97.977 ;
        RECT 0 91 5.5 98 ;
      LAYER MET3 ;
        RECT 0 91.983 6.5 97.017 ;
        RECT 0 91.943 6.466 97.057 ;
        RECT 0 91.897 6.42 97.103 ;
        RECT 0 91.851 6.374 97.149 ;
        RECT 0 91.805 6.328 97.195 ;
        RECT 0 91.759 6.282 97.241 ;
        RECT 0 91.713 6.236 97.287 ;
        RECT 0 91.667 6.19 97.333 ;
        RECT 0 91.621 6.144 97.379 ;
        RECT 0 91.575 6.098 97.425 ;
        RECT 0 91.529 6.052 97.471 ;
        RECT 0 91.483 6.006 97.517 ;
        RECT 0 91.437 5.96 97.563 ;
        RECT 0 91.391 5.914 97.609 ;
        RECT 0 91.345 5.868 97.655 ;
        RECT 0 91.299 5.822 97.701 ;
        RECT 0 91.253 5.776 97.747 ;
        RECT 0 91.207 5.73 97.793 ;
        RECT 0 91.161 5.684 97.839 ;
        RECT 0 91.115 5.638 97.885 ;
        RECT 0 91.069 5.592 97.931 ;
        RECT 0 91.023 5.546 97.977 ;
        RECT 0 91 5.5 98 ;
      LAYER MET2 ;
        RECT 0 91 65 98 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA2 ;
    ANTENNAPARTIALCUTAREA 1.539 LAYER VIA4 ;
    PORT
      LAYER MET5 ;
        RECT 0 78.5 65 89.5 ;
        RECT 0 3.788 1.5 15.212 ;
        RECT 0 3.753 1.476 15.247 ;
        RECT 0 3.707 1.43 15.293 ;
        RECT 0 3.661 1.384 15.339 ;
        RECT 0 3.615 1.338 15.385 ;
        RECT 0 3.569 1.292 15.431 ;
        RECT 0 3.523 1.246 15.477 ;
        RECT 0 3.5 1.2 15.5 ;
        RECT 0 17.288 1.5 28.712 ;
        RECT 0 17.253 1.476 28.747 ;
        RECT 0 17.207 1.43 28.793 ;
        RECT 0 17.161 1.384 28.839 ;
        RECT 0 17.115 1.338 28.885 ;
        RECT 0 17.069 1.292 28.931 ;
        RECT 0 17.023 1.246 28.977 ;
        RECT 0 17 1.2 29 ;
      LAYER MET4 ;
        RECT 0 79.483 6.5 88.517 ;
        RECT 0 79.443 6.466 88.557 ;
        RECT 0 79.397 6.42 88.603 ;
        RECT 0 79.351 6.374 88.649 ;
        RECT 0 79.305 6.328 88.695 ;
        RECT 0 79.259 6.282 88.741 ;
        RECT 0 79.213 6.236 88.787 ;
        RECT 0 79.167 6.19 88.833 ;
        RECT 0 79.121 6.144 88.879 ;
        RECT 0 79.075 6.098 88.925 ;
        RECT 0 79.029 6.052 88.971 ;
        RECT 0 78.983 6.006 89.017 ;
        RECT 0 78.937 5.96 89.063 ;
        RECT 0 78.891 5.914 89.109 ;
        RECT 0 78.845 5.868 89.155 ;
        RECT 0 78.799 5.822 89.201 ;
        RECT 0 78.753 5.776 89.247 ;
        RECT 0 78.707 5.73 89.293 ;
        RECT 0 78.661 5.684 89.339 ;
        RECT 0 78.615 5.638 89.385 ;
        RECT 0 78.569 5.592 89.431 ;
        RECT 0 78.523 5.546 89.477 ;
        RECT 0 78.5 5.5 89.5 ;
        RECT 0 3.788 1.5 15.212 ;
        RECT 0 3.753 1.476 15.247 ;
        RECT 0 3.707 1.43 15.293 ;
        RECT 0 3.661 1.384 15.339 ;
        RECT 0 3.615 1.338 15.385 ;
        RECT 0 3.569 1.292 15.431 ;
        RECT 0 3.523 1.246 15.477 ;
        RECT 0 3.5 1.2 15.5 ;
        RECT 0 17.288 1.5 28.712 ;
        RECT 0 17.253 1.476 28.747 ;
        RECT 0 17.207 1.43 28.793 ;
        RECT 0 17.161 1.384 28.839 ;
        RECT 0 17.115 1.338 28.885 ;
        RECT 0 17.069 1.292 28.931 ;
        RECT 0 17.023 1.246 28.977 ;
        RECT 0 17 1.2 29 ;
      LAYER MET3 ;
        RECT 0 79.483 6.5 88.517 ;
        RECT 0 79.443 6.466 88.557 ;
        RECT 0 79.397 6.42 88.603 ;
        RECT 0 79.351 6.374 88.649 ;
        RECT 0 79.305 6.328 88.695 ;
        RECT 0 79.259 6.282 88.741 ;
        RECT 0 79.213 6.236 88.787 ;
        RECT 0 79.167 6.19 88.833 ;
        RECT 0 79.121 6.144 88.879 ;
        RECT 0 79.075 6.098 88.925 ;
        RECT 0 79.029 6.052 88.971 ;
        RECT 0 78.983 6.006 89.017 ;
        RECT 0 78.937 5.96 89.063 ;
        RECT 0 78.891 5.914 89.109 ;
        RECT 0 78.845 5.868 89.155 ;
        RECT 0 78.799 5.822 89.201 ;
        RECT 0 78.753 5.776 89.247 ;
        RECT 0 78.707 5.73 89.293 ;
        RECT 0 78.661 5.684 89.339 ;
        RECT 0 78.615 5.638 89.385 ;
        RECT 0 78.569 5.592 89.431 ;
        RECT 0 78.523 5.546 89.477 ;
        RECT 0 78.5 5.5 89.5 ;
        RECT 0 3.788 1.5 15.212 ;
        RECT 0 3.753 1.476 15.247 ;
        RECT 0 3.707 1.43 15.293 ;
        RECT 0 3.661 1.384 15.339 ;
        RECT 0 3.615 1.338 15.385 ;
        RECT 0 3.569 1.292 15.431 ;
        RECT 0 3.523 1.246 15.477 ;
        RECT 0 3.5 1.2 15.5 ;
        RECT 0 17.288 1.5 28.712 ;
        RECT 0 17.253 1.476 28.747 ;
        RECT 0 17.207 1.43 28.793 ;
        RECT 0 17.161 1.384 28.839 ;
        RECT 0 17.115 1.338 28.885 ;
        RECT 0 17.069 1.292 28.931 ;
        RECT 0 17.023 1.246 28.977 ;
        RECT 0 17 1.2 29 ;
      LAYER MET2 ;
        RECT 0 17 65 29 ;
        RECT 0 3.5 65 15.5 ;
        RECT 59.805 3.5 60.995 29 ;
        RECT 54.225 3.5 55.415 29 ;
        RECT 48.645 3.5 49.835 29 ;
        RECT 43.065 3.5 44.255 29 ;
        RECT 37.485 3.5 38.675 29 ;
        RECT 31.905 3.5 33.095 29 ;
        RECT 26.325 3.5 27.515 29 ;
        RECT 20.745 3.5 21.935 29 ;
        RECT 15.165 3.5 16.355 29 ;
        RECT 9.585 3.5 10.775 29 ;
        RECT 4.005 3.5 5.195 29 ;
        RECT 0 78.5 65 89.5 ;
    END
  END VSSIO
  OBS
    LAYER MET1 SPACING 0.09 ;
      RECT 0 -20 65 110 ;
    LAYER MET2 SPACING 0.1 ;
      RECT 57.175 107.675 65 110 ;
      RECT 0 107.675 7.825 110 ;
      RECT 0 107.675 65 108.825 ;
      RECT 0 -20 65 3.325 ;
      RECT 61.17 15.675 65 16.825 ;
      RECT 0 29.175 65 30.325 ;
      RECT 59.38 42.675 65 43.825 ;
      RECT 59.38 56.175 65 57.325 ;
      RECT 0 63.675 65 68.325 ;
      RECT 0 77.175 65 78.325 ;
      RECT 0 89.675 65 90.825 ;
      RECT 0 98.175 65 99.325 ;
      RECT 55.59 15.675 59.63 16.825 ;
      RECT 53.8 42.675 55.84 43.825 ;
      RECT 53.8 56.175 55.84 57.325 ;
      RECT 50.01 15.675 54.05 16.825 ;
      RECT 48.22 42.675 50.26 43.825 ;
      RECT 48.22 56.175 50.26 57.325 ;
      RECT 44.43 15.675 48.47 16.825 ;
      RECT 42.64 42.675 44.68 43.825 ;
      RECT 42.64 56.175 44.68 57.325 ;
      RECT 38.85 15.675 42.89 16.825 ;
      RECT 37.06 42.675 39.1 43.825 ;
      RECT 37.06 56.175 39.1 57.325 ;
      RECT 33.27 15.675 37.31 16.825 ;
      RECT 31.48 42.675 33.52 43.825 ;
      RECT 31.48 56.175 33.52 57.325 ;
      RECT 27.69 15.675 31.73 16.825 ;
      RECT 25.9 42.675 27.94 43.825 ;
      RECT 25.9 56.175 27.94 57.325 ;
      RECT 22.11 15.675 26.15 16.825 ;
      RECT 20.32 42.675 22.36 43.825 ;
      RECT 20.32 56.175 22.36 57.325 ;
      RECT 16.53 15.675 20.57 16.825 ;
      RECT 14.74 42.675 16.78 43.825 ;
      RECT 14.74 56.175 16.78 57.325 ;
      RECT 10.95 15.675 14.99 16.825 ;
      RECT 9.16 42.675 11.2 43.825 ;
      RECT 9.16 56.175 11.2 57.325 ;
      RECT 5.37 15.675 9.41 16.825 ;
      RECT 0 42.675 5.62 43.825 ;
      RECT 0 56.175 5.62 57.325 ;
      RECT 0 15.675 3.83 16.825 ;
    LAYER MET3 SPACING 0.1 ;
      RECT 61.175 -20 65 3.335 ;
      RECT 1.375 -20 3.825 3.335 ;
      RECT 0 -20 3.825 3.325 ;
      RECT 0 -20 65 -0.175 ;
      RECT 63.8 3.5 65 15.5 ;
      RECT 63.776 3.512 65 15.488 ;
      RECT 63.73 3.547 65 15.453 ;
      RECT 63.684 3.593 65 15.407 ;
      RECT 63.638 3.639 65 15.361 ;
      RECT 63.592 3.685 65 15.315 ;
      RECT 63.546 3.731 65 15.269 ;
      RECT 63.5 3.777 65 15.223 ;
      RECT 63.8 17 65 29 ;
      RECT 63.776 17.012 65 28.988 ;
      RECT 63.73 17.047 65 28.953 ;
      RECT 63.684 17.093 65 28.907 ;
      RECT 63.638 17.139 65 28.861 ;
      RECT 63.592 17.185 65 28.815 ;
      RECT 63.546 17.231 65 28.769 ;
      RECT 63.5 17.277 65 28.723 ;
      RECT 59.466 78.517 59.5 89.483 ;
      RECT 59.42 78.557 59.466 89.443 ;
      RECT 59.374 78.603 59.42 89.397 ;
      RECT 59.328 78.649 59.374 89.351 ;
      RECT 59.282 78.695 59.328 89.305 ;
      RECT 59.236 78.741 59.282 89.259 ;
      RECT 59.19 78.787 59.236 89.213 ;
      RECT 59.144 78.833 59.19 89.167 ;
      RECT 59.098 78.879 59.144 89.121 ;
      RECT 59.052 78.925 59.098 89.075 ;
      RECT 59.006 78.971 59.052 89.029 ;
      RECT 58.96 79.017 59.006 88.983 ;
      RECT 58.914 79.063 58.96 88.937 ;
      RECT 58.868 79.109 58.914 88.891 ;
      RECT 58.822 79.155 58.868 88.845 ;
      RECT 58.776 79.201 58.822 88.799 ;
      RECT 58.73 79.247 58.776 88.753 ;
      RECT 58.684 79.293 58.73 88.707 ;
      RECT 58.638 79.339 58.684 88.661 ;
      RECT 58.592 79.385 58.638 88.615 ;
      RECT 58.546 79.431 58.592 88.569 ;
      RECT 58.5 79.477 58.546 88.523 ;
      RECT 59.5 78.5 65 89.5 ;
      RECT 59.466 91.017 59.5 97.983 ;
      RECT 59.42 91.057 59.466 97.943 ;
      RECT 59.374 91.103 59.42 97.897 ;
      RECT 59.328 91.149 59.374 97.851 ;
      RECT 59.282 91.195 59.328 97.805 ;
      RECT 59.236 91.241 59.282 97.759 ;
      RECT 59.19 91.287 59.236 97.713 ;
      RECT 59.144 91.333 59.19 97.667 ;
      RECT 59.098 91.379 59.144 97.621 ;
      RECT 59.052 91.425 59.098 97.575 ;
      RECT 59.006 91.471 59.052 97.529 ;
      RECT 58.96 91.517 59.006 97.483 ;
      RECT 58.914 91.563 58.96 97.437 ;
      RECT 58.868 91.609 58.914 97.391 ;
      RECT 58.822 91.655 58.868 97.345 ;
      RECT 58.776 91.701 58.822 97.299 ;
      RECT 58.73 91.747 58.776 97.253 ;
      RECT 58.684 91.793 58.73 97.207 ;
      RECT 58.638 91.839 58.684 97.161 ;
      RECT 58.592 91.885 58.638 97.115 ;
      RECT 58.546 91.931 58.592 97.069 ;
      RECT 58.5 91.977 58.546 97.023 ;
      RECT 59.5 91 65 98 ;
      RECT 59.466 99.517 59.5 107.483 ;
      RECT 59.42 99.557 59.466 107.443 ;
      RECT 59.374 99.603 59.42 107.397 ;
      RECT 59.328 99.649 59.374 107.351 ;
      RECT 59.282 99.695 59.328 107.305 ;
      RECT 59.236 99.741 59.282 107.259 ;
      RECT 59.19 99.787 59.236 107.213 ;
      RECT 59.144 99.833 59.19 107.167 ;
      RECT 59.098 99.879 59.144 107.121 ;
      RECT 59.052 99.925 59.098 107.075 ;
      RECT 59.006 99.971 59.052 107.029 ;
      RECT 58.96 100.017 59.006 106.983 ;
      RECT 58.914 100.063 58.96 106.937 ;
      RECT 58.868 100.109 58.914 106.891 ;
      RECT 58.822 100.155 58.868 106.845 ;
      RECT 58.776 100.201 58.822 106.799 ;
      RECT 58.73 100.247 58.776 106.753 ;
      RECT 58.684 100.293 58.73 106.707 ;
      RECT 58.638 100.339 58.684 106.661 ;
      RECT 58.592 100.385 58.638 106.615 ;
      RECT 58.546 100.431 58.592 106.569 ;
      RECT 58.5 100.477 58.546 106.523 ;
      RECT 59.5 99.5 65 107.5 ;
      RECT 5.675 77.175 7.825 78.335 ;
      RECT 0 77.175 7.825 78.325 ;
      RECT 5.675 89.665 7.825 90.835 ;
      RECT 0 89.675 7.825 90.825 ;
      RECT 5.675 98.165 7.825 99.335 ;
      RECT 0 98.175 7.825 99.325 ;
      RECT 0 107.675 7.825 110 ;
      RECT 5.675 107.665 7.825 110 ;
      RECT 1.375 15.665 2.825 16.835 ;
      RECT 0 15.675 2.825 16.825 ;
      RECT 0 29.175 2.825 30.325 ;
      RECT 1.375 29.165 2.825 30.325 ;
      RECT 62.175 15.665 65 16.835 ;
      RECT 62.175 29.165 65 30.325 ;
      RECT 62.175 42.675 65 43.825 ;
      RECT 62.175 56.175 65 57.325 ;
      RECT 58.175 63.675 65 68.325 ;
      RECT 57.175 77.175 65 78.335 ;
      RECT 57.175 89.665 65 90.835 ;
      RECT 57.175 98.165 65 99.335 ;
      RECT 57.175 107.665 65 110 ;
      RECT 55.58 15.665 56.825 16.835 ;
      RECT 50.675 29.165 56.825 30.335 ;
      RECT 53.79 42.665 55.85 43.835 ;
      RECT 53.79 56.165 55.85 57.335 ;
      RECT 50.675 15.665 54.06 16.835 ;
      RECT 44.515 63.675 45.825 68.325 ;
      RECT 44.515 77.175 45.825 78.335 ;
      RECT 44.515 89.665 45.825 90.835 ;
      RECT 44.515 98.165 45.825 99.335 ;
      RECT 44.515 107.665 45.825 108.825 ;
      RECT 38.84 15.665 42.825 16.835 ;
      RECT 36.675 29.165 42.825 30.335 ;
      RECT 42.63 42.665 42.825 43.835 ;
      RECT 42.63 56.165 42.825 57.335 ;
      RECT 37.05 42.665 39.11 43.835 ;
      RECT 37.05 56.165 39.11 57.335 ;
      RECT 36.675 15.665 37.32 16.835 ;
      RECT 31.835 63.675 33.095 68.325 ;
      RECT 31.835 77.175 33.095 78.335 ;
      RECT 31.835 89.665 33.095 90.835 ;
      RECT 31.835 98.165 33.095 99.335 ;
      RECT 31.835 107.665 33.095 108.825 ;
      RECT 27.68 15.665 28.825 16.835 ;
      RECT 22.675 29.165 28.825 30.335 ;
      RECT 25.89 42.665 27.95 43.835 ;
      RECT 25.89 56.165 27.95 57.335 ;
      RECT 22.675 15.665 26.16 16.835 ;
      RECT 19.175 63.675 20.485 68.325 ;
      RECT 19.175 77.175 20.485 78.335 ;
      RECT 19.175 89.665 20.485 90.835 ;
      RECT 19.175 98.165 20.485 99.335 ;
      RECT 19.175 107.665 20.485 108.825 ;
      RECT 10.94 15.665 14.825 16.835 ;
      RECT 8.675 29.165 14.825 30.335 ;
      RECT 9.15 42.665 11.21 43.835 ;
      RECT 9.15 56.165 11.21 57.335 ;
      RECT 8.675 15.665 9.42 16.835 ;
      RECT 0 63.675 6.825 68.325 ;
      RECT 0 42.675 2.825 43.825 ;
      RECT 0 56.175 2.825 57.325 ;
    LAYER MET4 SPACING 0.1 ;
      RECT 62.175 -20 65 30.325 ;
      RECT 0 29.175 2.825 30.325 ;
      RECT 1.675 -20 2.825 30.325 ;
      RECT 1.375 29.152 2.825 30.325 ;
      RECT 1.651 28.887 2.825 30.325 ;
      RECT 1.421 29.106 2.825 30.325 ;
      RECT 1.605 28.922 2.825 30.325 ;
      RECT 1.467 29.06 2.825 30.325 ;
      RECT 1.559 28.968 2.825 30.325 ;
      RECT 1.513 29.014 2.825 30.325 ;
      RECT 1.651 15.387 2.825 17.113 ;
      RECT 1.605 15.422 2.825 17.078 ;
      RECT 1.559 15.468 2.825 17.032 ;
      RECT 1.513 15.514 2.825 16.986 ;
      RECT 1.467 15.56 2.825 16.94 ;
      RECT 1.421 15.606 2.825 16.894 ;
      RECT 1.375 15.652 2.825 16.848 ;
      RECT 0 15.675 2.825 16.825 ;
      RECT 62.141 -20 65 4.308 ;
      RECT 1.675 -20 2.871 4.302 ;
      RECT 62.095 -20 65 4.268 ;
      RECT 1.675 -20 2.917 4.256 ;
      RECT 62.049 -20 65 4.222 ;
      RECT 1.675 -20 2.963 4.21 ;
      RECT 62.003 -20 65 4.176 ;
      RECT 1.675 -20 3.009 4.164 ;
      RECT 61.957 -20 65 4.13 ;
      RECT 1.675 -20 3.055 4.118 ;
      RECT 61.911 -20 65 4.084 ;
      RECT 1.675 -20 3.101 4.072 ;
      RECT 61.865 -20 65 4.038 ;
      RECT 1.675 -20 3.147 4.026 ;
      RECT 61.819 -20 65 3.992 ;
      RECT 1.675 -20 3.193 3.98 ;
      RECT 61.773 -20 65 3.946 ;
      RECT 1.675 -20 3.239 3.934 ;
      RECT 61.727 -20 65 3.9 ;
      RECT 1.675 -20 3.285 3.888 ;
      RECT 61.681 -20 65 3.854 ;
      RECT 1.675 -20 3.331 3.842 ;
      RECT 61.635 -20 65 3.808 ;
      RECT 1.675 -20 3.377 3.796 ;
      RECT 61.589 -20 65 3.762 ;
      RECT 1.675 -20 3.423 3.75 ;
      RECT 61.543 -20 65 3.716 ;
      RECT 1.675 -20 3.469 3.704 ;
      RECT 61.497 -20 65 3.67 ;
      RECT 1.675 -20 3.515 3.658 ;
      RECT 61.451 -20 65 3.624 ;
      RECT 1.651 -20 3.515 3.613 ;
      RECT 1.651 -20 3.561 3.612 ;
      RECT 61.405 -20 65 3.578 ;
      RECT 1.605 -20 3.561 3.578 ;
      RECT 1.605 -20 3.607 3.566 ;
      RECT 61.359 -20 65 3.532 ;
      RECT 1.559 -20 3.607 3.532 ;
      RECT 1.559 -20 3.653 3.52 ;
      RECT 61.313 -20 65 3.486 ;
      RECT 1.513 -20 3.653 3.486 ;
      RECT 1.513 -20 3.699 3.474 ;
      RECT 61.267 -20 65 3.44 ;
      RECT 1.467 -20 3.699 3.44 ;
      RECT 1.467 -20 3.745 3.428 ;
      RECT 61.221 -20 65 3.394 ;
      RECT 1.421 -20 3.745 3.394 ;
      RECT 1.421 -20 3.791 3.382 ;
      RECT 61.175 -20 65 3.348 ;
      RECT 1.375 -20 3.791 3.348 ;
      RECT 1.375 -20 3.825 3.342 ;
      RECT 0 -20 3.825 3.325 ;
      RECT 0 -20 65 -0.175 ;
      RECT 0 107.675 7.825 110 ;
      RECT 6.675 77.175 7.825 110 ;
      RECT 5.675 107.652 7.825 110 ;
      RECT 6.641 106.692 7.825 110 ;
      RECT 5.721 107.606 7.825 110 ;
      RECT 6.595 106.732 7.825 110 ;
      RECT 5.767 107.56 7.825 110 ;
      RECT 6.549 106.778 7.825 110 ;
      RECT 5.813 107.514 7.825 110 ;
      RECT 6.503 106.824 7.825 110 ;
      RECT 5.859 107.468 7.825 110 ;
      RECT 6.457 106.87 7.825 110 ;
      RECT 5.905 107.422 7.825 110 ;
      RECT 6.411 106.916 7.825 110 ;
      RECT 5.951 107.376 7.825 110 ;
      RECT 6.365 106.962 7.825 110 ;
      RECT 5.997 107.33 7.825 110 ;
      RECT 6.319 107.008 7.825 110 ;
      RECT 6.043 107.284 7.825 110 ;
      RECT 6.273 107.054 7.825 110 ;
      RECT 6.089 107.238 7.825 110 ;
      RECT 6.227 107.1 7.825 110 ;
      RECT 6.135 107.192 7.825 110 ;
      RECT 6.181 107.146 7.825 110 ;
      RECT 6.641 97.192 7.825 100.308 ;
      RECT 6.595 97.232 7.825 100.268 ;
      RECT 6.549 97.278 7.825 100.222 ;
      RECT 6.503 97.324 7.825 100.176 ;
      RECT 6.457 97.37 7.825 100.13 ;
      RECT 6.411 97.416 7.825 100.084 ;
      RECT 6.365 97.462 7.825 100.038 ;
      RECT 6.319 97.508 7.825 99.992 ;
      RECT 6.273 97.554 7.825 99.946 ;
      RECT 6.227 97.6 7.825 99.9 ;
      RECT 6.181 97.646 7.825 99.854 ;
      RECT 6.135 97.692 7.825 99.808 ;
      RECT 6.089 97.738 7.825 99.762 ;
      RECT 6.043 97.784 7.825 99.716 ;
      RECT 5.997 97.83 7.825 99.67 ;
      RECT 5.951 97.876 7.825 99.624 ;
      RECT 5.905 97.922 7.825 99.578 ;
      RECT 5.859 97.968 7.825 99.532 ;
      RECT 5.813 98.014 7.825 99.486 ;
      RECT 5.767 98.06 7.825 99.44 ;
      RECT 5.721 98.106 7.825 99.394 ;
      RECT 5.675 98.152 7.825 99.348 ;
      RECT 0 98.175 7.825 99.325 ;
      RECT 6.641 88.692 7.825 91.808 ;
      RECT 6.595 88.732 7.825 91.768 ;
      RECT 6.549 88.778 7.825 91.722 ;
      RECT 6.503 88.824 7.825 91.676 ;
      RECT 6.457 88.87 7.825 91.63 ;
      RECT 6.411 88.916 7.825 91.584 ;
      RECT 6.365 88.962 7.825 91.538 ;
      RECT 6.319 89.008 7.825 91.492 ;
      RECT 6.273 89.054 7.825 91.446 ;
      RECT 6.227 89.1 7.825 91.4 ;
      RECT 6.181 89.146 7.825 91.354 ;
      RECT 6.135 89.192 7.825 91.308 ;
      RECT 6.089 89.238 7.825 91.262 ;
      RECT 6.043 89.284 7.825 91.216 ;
      RECT 5.997 89.33 7.825 91.17 ;
      RECT 5.951 89.376 7.825 91.124 ;
      RECT 5.905 89.422 7.825 91.078 ;
      RECT 5.859 89.468 7.825 91.032 ;
      RECT 5.813 89.514 7.825 90.986 ;
      RECT 5.767 89.56 7.825 90.94 ;
      RECT 5.721 89.606 7.825 90.894 ;
      RECT 5.675 89.652 7.825 90.848 ;
      RECT 0 89.675 7.825 90.825 ;
      RECT 6.641 77.175 7.825 79.308 ;
      RECT 6.595 77.175 7.825 79.268 ;
      RECT 6.549 77.175 7.825 79.222 ;
      RECT 6.503 77.175 7.825 79.176 ;
      RECT 6.457 77.175 7.825 79.13 ;
      RECT 6.411 77.175 7.825 79.084 ;
      RECT 6.365 77.175 7.825 79.038 ;
      RECT 6.319 77.175 7.825 78.992 ;
      RECT 6.273 77.175 7.825 78.946 ;
      RECT 6.227 77.175 7.825 78.9 ;
      RECT 6.181 77.175 7.825 78.854 ;
      RECT 6.135 77.175 7.825 78.808 ;
      RECT 6.089 77.175 7.825 78.762 ;
      RECT 6.043 77.175 7.825 78.716 ;
      RECT 5.997 77.175 7.825 78.67 ;
      RECT 5.951 77.175 7.825 78.624 ;
      RECT 5.905 77.175 7.825 78.578 ;
      RECT 5.859 77.175 7.825 78.532 ;
      RECT 5.813 77.175 7.825 78.486 ;
      RECT 5.767 77.175 7.825 78.44 ;
      RECT 5.721 77.175 7.825 78.394 ;
      RECT 5.675 77.175 7.825 78.348 ;
      RECT 0 77.175 7.825 78.325 ;
      RECT 62.175 42.675 65 43.825 ;
      RECT 62.175 56.175 65 57.325 ;
      RECT 58.175 63.675 65 68.325 ;
      RECT 57.175 77.175 65 110 ;
      RECT 50.675 12.175 56.825 18.905 ;
      RECT 50.675 26.755 56.825 32.905 ;
      RECT 50.675 40.755 56.825 46.905 ;
      RECT 50.675 54.755 56.825 60.905 ;
      RECT 44.515 63.675 45.825 68.325 ;
      RECT 44.515 77.175 45.825 108.825 ;
      RECT 36.675 12.175 42.825 18.905 ;
      RECT 36.675 26.755 42.825 32.905 ;
      RECT 36.675 40.755 42.825 46.905 ;
      RECT 36.675 54.755 42.825 60.905 ;
      RECT 31.835 63.675 33.095 68.325 ;
      RECT 31.835 77.175 33.095 108.825 ;
      RECT 22.675 12.175 28.825 18.905 ;
      RECT 22.675 26.755 28.825 32.905 ;
      RECT 22.675 40.755 28.825 46.905 ;
      RECT 22.675 54.755 28.825 60.905 ;
      RECT 19.175 63.675 20.485 68.325 ;
      RECT 19.175 77.175 20.485 108.825 ;
      RECT 8.675 12.175 14.825 18.905 ;
      RECT 8.675 26.755 14.825 32.905 ;
      RECT 8.675 40.755 14.825 46.905 ;
      RECT 8.675 54.755 14.825 60.905 ;
      RECT 0 63.675 6.825 68.325 ;
      RECT 0 42.675 2.825 43.825 ;
      RECT 0 56.175 2.825 57.325 ;
    LAYER MET5 SPACING 0.1 ;
      RECT 62.33 -20 65 30.17 ;
      RECT 0 29.33 2.67 30.17 ;
      RECT 1.83 -20 2.67 30.17 ;
      RECT 1.53 29.307 2.67 30.17 ;
      RECT 1.806 29.042 2.67 30.17 ;
      RECT 1.576 29.261 2.67 30.17 ;
      RECT 1.76 29.077 2.67 30.17 ;
      RECT 1.622 29.215 2.67 30.17 ;
      RECT 1.714 29.123 2.67 30.17 ;
      RECT 1.668 29.169 2.67 30.17 ;
      RECT 1.806 15.542 2.67 16.958 ;
      RECT 1.76 15.577 2.67 16.923 ;
      RECT 1.714 15.623 2.67 16.877 ;
      RECT 1.668 15.669 2.67 16.831 ;
      RECT 1.622 15.715 2.67 16.785 ;
      RECT 1.576 15.761 2.67 16.739 ;
      RECT 1.53 15.807 2.67 16.693 ;
      RECT 0 15.83 2.67 16.67 ;
      RECT 62.296 -20 65 4.153 ;
      RECT 1.83 -20 2.716 4.147 ;
      RECT 62.25 -20 65 4.113 ;
      RECT 1.83 -20 2.762 4.101 ;
      RECT 62.204 -20 65 4.067 ;
      RECT 1.83 -20 2.808 4.055 ;
      RECT 62.158 -20 65 4.021 ;
      RECT 1.83 -20 2.854 4.009 ;
      RECT 62.112 -20 65 3.975 ;
      RECT 1.83 -20 2.9 3.963 ;
      RECT 62.066 -20 65 3.929 ;
      RECT 1.83 -20 2.946 3.917 ;
      RECT 62.02 -20 65 3.883 ;
      RECT 1.83 -20 2.992 3.871 ;
      RECT 61.974 -20 65 3.837 ;
      RECT 1.83 -20 3.038 3.825 ;
      RECT 61.928 -20 65 3.791 ;
      RECT 1.83 -20 3.084 3.779 ;
      RECT 61.882 -20 65 3.745 ;
      RECT 1.83 -20 3.13 3.733 ;
      RECT 61.836 -20 65 3.699 ;
      RECT 1.83 -20 3.176 3.687 ;
      RECT 61.79 -20 65 3.653 ;
      RECT 1.83 -20 3.222 3.641 ;
      RECT 61.744 -20 65 3.607 ;
      RECT 1.83 -20 3.268 3.595 ;
      RECT 61.698 -20 65 3.561 ;
      RECT 1.83 -20 3.314 3.549 ;
      RECT 61.652 -20 65 3.515 ;
      RECT 1.83 -20 3.36 3.503 ;
      RECT 61.606 -20 65 3.469 ;
      RECT 1.806 -20 3.36 3.458 ;
      RECT 1.806 -20 3.406 3.457 ;
      RECT 61.56 -20 65 3.423 ;
      RECT 1.76 -20 3.406 3.423 ;
      RECT 1.76 -20 3.452 3.411 ;
      RECT 61.514 -20 65 3.377 ;
      RECT 1.714 -20 3.452 3.377 ;
      RECT 1.714 -20 3.498 3.365 ;
      RECT 61.468 -20 65 3.331 ;
      RECT 1.668 -20 3.498 3.331 ;
      RECT 1.668 -20 3.544 3.319 ;
      RECT 61.422 -20 65 3.285 ;
      RECT 1.622 -20 3.544 3.285 ;
      RECT 1.622 -20 3.59 3.273 ;
      RECT 61.376 -20 65 3.239 ;
      RECT 1.576 -20 3.59 3.239 ;
      RECT 1.576 -20 3.636 3.227 ;
      RECT 61.33 -20 65 3.193 ;
      RECT 1.53 -20 3.636 3.193 ;
      RECT 1.53 -20 3.67 3.187 ;
      RECT 0 -20 3.67 3.17 ;
      RECT 0 -20 65 -0.33 ;
      RECT 57.33 107.83 65 110 ;
      RECT 57.165 107.83 65 108.67 ;
      RECT 0 107.83 7.67 110 ;
      RECT 0 107.83 7.835 108.67 ;
      RECT 62.33 42.83 65 43.67 ;
      RECT 62.33 56.33 65 57.17 ;
      RECT 58.33 63.83 65 68.17 ;
      RECT 57.165 77.33 65 78.17 ;
      RECT 57.165 89.83 65 90.67 ;
      RECT 57.165 98.33 65 99.17 ;
      RECT 50.83 12.33 56.67 18.75 ;
      RECT 50.83 26.91 56.67 32.75 ;
      RECT 50.83 40.91 56.67 46.75 ;
      RECT 50.83 54.91 56.67 60.75 ;
      RECT 44.505 77.33 45.835 78.17 ;
      RECT 44.505 89.83 45.835 90.67 ;
      RECT 44.505 98.33 45.835 99.17 ;
      RECT 44.505 107.83 45.835 108.67 ;
      RECT 44.67 63.83 45.67 68.17 ;
      RECT 36.83 12.33 42.67 18.75 ;
      RECT 36.83 26.91 42.67 32.75 ;
      RECT 36.83 40.91 42.67 46.75 ;
      RECT 36.83 54.91 42.67 60.75 ;
      RECT 31.825 77.33 33.105 78.17 ;
      RECT 31.825 89.83 33.105 90.67 ;
      RECT 31.825 98.33 33.105 99.17 ;
      RECT 31.825 107.83 33.105 108.67 ;
      RECT 31.99 63.83 32.94 68.17 ;
      RECT 22.83 12.33 28.67 18.75 ;
      RECT 22.83 26.91 28.67 32.75 ;
      RECT 22.83 40.91 28.67 46.75 ;
      RECT 22.83 54.91 28.67 60.75 ;
      RECT 19.165 77.33 20.495 78.17 ;
      RECT 19.165 89.83 20.495 90.67 ;
      RECT 19.165 98.33 20.495 99.17 ;
      RECT 19.165 107.83 20.495 108.67 ;
      RECT 19.33 63.83 20.33 68.17 ;
      RECT 8.83 12.33 14.67 18.75 ;
      RECT 8.83 26.91 14.67 32.75 ;
      RECT 8.83 40.91 14.67 46.75 ;
      RECT 8.83 54.91 14.67 60.75 ;
      RECT 0 77.33 7.835 78.17 ;
      RECT 0 89.83 7.835 90.67 ;
      RECT 0 98.33 7.835 99.17 ;
      RECT 0 63.83 6.67 68.17 ;
      RECT 0 42.83 2.67 43.67 ;
      RECT 0 56.33 2.67 57.17 ;
    LAYER T4M2 SPACING 0.4 ;
      RECT 64.576 -20 65 0.444 ;
      RECT 0 -20 0.436 0.427 ;
      RECT 64.53 -20 65 0.398 ;
      RECT 0 -20 0.482 0.381 ;
      RECT 64.484 -20 65 0.352 ;
      RECT 0 -20 0.528 0.335 ;
      RECT 64.438 -20 65 0.306 ;
      RECT 0 -20 0.574 0.289 ;
      RECT 64.392 -20 65 0.26 ;
      RECT 0 -20 0.62 0.243 ;
      RECT 64.346 -20 65 0.214 ;
      RECT 0 -20 0.666 0.197 ;
      RECT 64.3 -20 65 0.168 ;
      RECT 0 -20 0.7 0.157 ;
      RECT 0 -20 65 -3.3 ;
      RECT 57.6 108.1 65 110 ;
      RECT 0 108.1 7.4 110 ;
    LAYER RDL SPACING 2 ;
      RECT 0 -20 65 -4.9 ;
      RECT 0 81.9 65 110 ;
      RECT 3 4.5 62 63.5 ;
  END
END P65_1233_VDDIO3

MACRO P65_1233_VSS1
  CLASS PAD ;
  ORIGIN 0 20 ;
  FOREIGN P65_1233_VSS1 0 -20 ;
  SIZE 65 BY 130 ;
  SYMMETRY X Y R90 ;
  SITE IOSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER MET5 ;
        RECT 0 99.5 65 107.5 ;
      LAYER MET4 ;
        RECT 0 99.5 65 107.5 ;
      LAYER MET3 ;
        RECT 0 99.5 65 107.5 ;
      LAYER MET2 ;
        RECT 0 99.5 65 107.5 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET5 ;
        RECT 0 68.5 65 77 ;
        RECT 0 30.788 1.5 42.212 ;
        RECT 0 30.753 1.476 42.247 ;
        RECT 0 30.707 1.43 42.293 ;
        RECT 0 30.661 1.384 42.339 ;
        RECT 0 30.615 1.338 42.385 ;
        RECT 0 30.569 1.292 42.431 ;
        RECT 0 30.523 1.246 42.477 ;
        RECT 0 30.5 1.2 42.5 ;
        RECT 0 44.288 1.5 55.712 ;
        RECT 0 44.253 1.476 55.747 ;
        RECT 0 44.207 1.43 55.793 ;
        RECT 0 44.161 1.384 55.839 ;
        RECT 0 44.115 1.338 55.885 ;
        RECT 0 44.069 1.292 55.931 ;
        RECT 0 44.023 1.246 55.977 ;
        RECT 0 44 1.2 56 ;
        RECT 0 57.788 1.5 63.212 ;
        RECT 0 57.753 1.476 63.247 ;
        RECT 0 57.707 1.43 63.293 ;
        RECT 0 57.661 1.384 63.339 ;
        RECT 0 57.615 1.338 63.385 ;
        RECT 0 57.569 1.292 63.431 ;
        RECT 0 57.523 1.246 63.477 ;
        RECT 0 57.5 1.2 63.5 ;
      LAYER MET4 ;
        RECT 0 68.5 65 77 ;
        RECT 0 30.788 1.5 42.212 ;
        RECT 0 30.753 1.476 42.247 ;
        RECT 0 30.707 1.43 42.293 ;
        RECT 0 30.661 1.384 42.339 ;
        RECT 0 30.615 1.338 42.385 ;
        RECT 0 30.569 1.292 42.431 ;
        RECT 0 30.523 1.246 42.477 ;
        RECT 0 30.5 1.2 42.5 ;
        RECT 0 44.288 1.5 55.712 ;
        RECT 0 44.253 1.476 55.747 ;
        RECT 0 44.207 1.43 55.793 ;
        RECT 0 44.161 1.384 55.839 ;
        RECT 0 44.115 1.338 55.885 ;
        RECT 0 44.069 1.292 55.931 ;
        RECT 0 44.023 1.246 55.977 ;
        RECT 0 44 1.2 56 ;
        RECT 0 57.788 1.5 63.212 ;
        RECT 0 57.753 1.476 63.247 ;
        RECT 0 57.707 1.43 63.293 ;
        RECT 0 57.661 1.384 63.339 ;
        RECT 0 57.615 1.338 63.385 ;
        RECT 0 57.569 1.292 63.431 ;
        RECT 0 57.523 1.246 63.477 ;
        RECT 0 57.5 1.2 63.5 ;
      LAYER MET3 ;
        RECT 0 68.5 65 77 ;
        RECT 0 30.788 1.5 42.212 ;
        RECT 0 30.753 1.476 42.247 ;
        RECT 0 30.707 1.43 42.293 ;
        RECT 0 30.661 1.384 42.339 ;
        RECT 0 30.615 1.338 42.385 ;
        RECT 0 30.569 1.292 42.431 ;
        RECT 0 30.523 1.246 42.477 ;
        RECT 0 30.5 1.2 42.5 ;
        RECT 0 44.288 1.5 55.712 ;
        RECT 0 44.253 1.476 55.747 ;
        RECT 0 44.207 1.43 55.793 ;
        RECT 0 44.161 1.384 55.839 ;
        RECT 0 44.115 1.338 55.885 ;
        RECT 0 44.069 1.292 55.931 ;
        RECT 0 44.023 1.246 55.977 ;
        RECT 0 44 1.2 56 ;
        RECT 0 57.788 1.5 63.212 ;
        RECT 0 57.753 1.476 63.247 ;
        RECT 0 57.707 1.43 63.293 ;
        RECT 0 57.661 1.384 63.339 ;
        RECT 0 57.615 1.338 63.385 ;
        RECT 0 57.569 1.292 63.431 ;
        RECT 0 57.523 1.246 63.477 ;
        RECT 0 57.5 1.2 63.5 ;
      LAYER MET2 ;
        RECT 0 57.5 65 63.5 ;
        RECT 0 44 65 56 ;
        RECT 0 30.5 65 42.5 ;
        RECT 54.5 30.5 56.5 63.5 ;
        RECT 49.9 30.5 51.9 63.5 ;
        RECT 45.3 30.5 47.3 63.5 ;
        RECT 40.7 30.5 42.7 63.5 ;
        RECT 36.1 30.5 38.1 63.5 ;
        RECT 31.5 30.5 33.5 63.5 ;
        RECT 26.9 30.5 28.9 63.5 ;
        RECT 22.3 30.5 24.3 63.5 ;
        RECT 17.7 30.5 19.7 63.5 ;
        RECT 13.1 30.5 15.1 63.5 ;
        RECT 8.5 30.5 10.5 63.5 ;
        RECT 0 68.5 65 77 ;
    END
  END VDDIO
  PIN VSS
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 6.2694 LAYER VIA4 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 5.1192 LAYER VIA2 ;
    PORT
      LAYER MET5 ;
        RECT 0 91 65 98 ;
      LAYER MET4 ;
        RECT 0 91 65 98 ;
      LAYER MET3 ;
        RECT 0 91 65 98 ;
      LAYER MET2 ;
        RECT 0 91 65 98 ;
    END
  END VSS
  PIN VSS1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3275 LAYER MET3 ;
    ANTENNAPARTIALMETALAREA 118 LAYER MET2 ;
    ANTENNAPARTIALMETALAREA 3275 LAYER MET4 ;
    ANTENNAPARTIALMETALAREA 3275 LAYER MET5 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA2 ;
    ANTENNAPARTIALCUTAREA 3.6207 LAYER VIA4 ;
    ANTENNAPARTIALCUTAREA 34.2144 LAYER T4V2 ;
    PORT
      LAYER T4M2 ;
        RECT 57 0.983 62 66.017 ;
        RECT 57 0.943 61.966 66.057 ;
        RECT 57 0.897 61.92 66.103 ;
        RECT 57 0.851 61.874 66.149 ;
        RECT 57 0.805 61.828 66.195 ;
        RECT 57 0.759 61.782 66.241 ;
        RECT 57 0.713 61.736 66.287 ;
        RECT 57 0.667 61.69 66.333 ;
        RECT 57 0.621 61.644 66.379 ;
        RECT 57 0.575 61.598 66.425 ;
        RECT 57 0.529 61.552 66.471 ;
        RECT 57 0.483 61.506 66.517 ;
        RECT 57 0.437 61.46 66.563 ;
        RECT 57 0.391 61.414 66.609 ;
        RECT 57 0.345 61.368 66.655 ;
        RECT 57 0.299 61.322 66.701 ;
        RECT 57 0.253 61.276 66.747 ;
        RECT 57 0.207 61.23 66.793 ;
        RECT 57 0.161 61.184 66.839 ;
        RECT 57 0.115 61.138 66.885 ;
        RECT 57 0.069 61.092 66.931 ;
        RECT 57 0.023 61.046 66.977 ;
        RECT 4 57.5 61 67 ;
        RECT 3 43.5 62 51 ;
        RECT 3 29.5 62 37 ;
        RECT 3 15.5 62 23 ;
        RECT 4 0 61 9 ;
        RECT 43 0 50.5 67 ;
        RECT 29 0 36.5 67 ;
        RECT 15 0 22.5 67 ;
        RECT 3 0.977 8.5 66.023 ;
        RECT 3.966 0.017 8.5 66.983 ;
        RECT 3.92 0.057 8.5 66.943 ;
        RECT 3.874 0.103 8.5 66.897 ;
        RECT 3.828 0.149 8.5 66.851 ;
        RECT 3.782 0.195 8.5 66.805 ;
        RECT 3.736 0.241 8.5 66.759 ;
        RECT 3.69 0.287 8.5 66.713 ;
        RECT 3.644 0.333 8.5 66.667 ;
        RECT 3.598 0.379 8.5 66.621 ;
        RECT 3.552 0.425 8.5 66.575 ;
        RECT 3.506 0.471 8.5 66.529 ;
        RECT 3.46 0.517 8.5 66.483 ;
        RECT 3.414 0.563 8.5 66.437 ;
        RECT 3.368 0.609 8.5 66.391 ;
        RECT 3.322 0.655 8.5 66.345 ;
        RECT 3.276 0.701 8.5 66.299 ;
        RECT 3.23 0.747 8.5 66.253 ;
        RECT 3.184 0.793 8.5 66.207 ;
        RECT 3.138 0.839 8.5 66.161 ;
        RECT 3.092 0.885 8.5 66.115 ;
        RECT 3.046 0.931 8.5 66.069 ;
      LAYER MET5 ;
        RECT 6.7 109 58.3 110 ;
      LAYER MET4 ;
        RECT 6.7 109 58.3 110 ;
      LAYER MET3 ;
        RECT 6.7 109 58.3 110 ;
      LAYER MET2 ;
        RECT 6.7 109 58.3 110 ;
    END
  END VSS1
  PIN VSSIO
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA2 ;
    ANTENNAPARTIALCUTAREA 9.7524 LAYER VIA4 ;
    PORT
      LAYER MET5 ;
        RECT 0 78.5 65 89.5 ;
        RECT 0 3.788 1.5 15.212 ;
        RECT 0 3.753 1.476 15.247 ;
        RECT 0 3.707 1.43 15.293 ;
        RECT 0 3.661 1.384 15.339 ;
        RECT 0 3.615 1.338 15.385 ;
        RECT 0 3.569 1.292 15.431 ;
        RECT 0 3.523 1.246 15.477 ;
        RECT 0 3.5 1.2 15.5 ;
        RECT 0 17.288 1.5 28.712 ;
        RECT 0 17.253 1.476 28.747 ;
        RECT 0 17.207 1.43 28.793 ;
        RECT 0 17.161 1.384 28.839 ;
        RECT 0 17.115 1.338 28.885 ;
        RECT 0 17.069 1.292 28.931 ;
        RECT 0 17.023 1.246 28.977 ;
        RECT 0 17 1.2 29 ;
      LAYER MET4 ;
        RECT 0 78.5 65 89.5 ;
        RECT 0 3.788 1.5 15.212 ;
        RECT 0 3.753 1.476 15.247 ;
        RECT 0 3.707 1.43 15.293 ;
        RECT 0 3.661 1.384 15.339 ;
        RECT 0 3.615 1.338 15.385 ;
        RECT 0 3.569 1.292 15.431 ;
        RECT 0 3.523 1.246 15.477 ;
        RECT 0 3.5 1.2 15.5 ;
        RECT 0 17.288 1.5 28.712 ;
        RECT 0 17.253 1.476 28.747 ;
        RECT 0 17.207 1.43 28.793 ;
        RECT 0 17.161 1.384 28.839 ;
        RECT 0 17.115 1.338 28.885 ;
        RECT 0 17.069 1.292 28.931 ;
        RECT 0 17.023 1.246 28.977 ;
        RECT 0 17 1.2 29 ;
      LAYER MET3 ;
        RECT 0 78.5 65 89.5 ;
        RECT 0 3.788 1.5 15.212 ;
        RECT 0 3.753 1.476 15.247 ;
        RECT 0 3.707 1.43 15.293 ;
        RECT 0 3.661 1.384 15.339 ;
        RECT 0 3.615 1.338 15.385 ;
        RECT 0 3.569 1.292 15.431 ;
        RECT 0 3.523 1.246 15.477 ;
        RECT 0 3.5 1.2 15.5 ;
        RECT 0 17.288 1.5 28.712 ;
        RECT 0 17.253 1.476 28.747 ;
        RECT 0 17.207 1.43 28.793 ;
        RECT 0 17.161 1.384 28.839 ;
        RECT 0 17.115 1.338 28.885 ;
        RECT 0 17.069 1.292 28.931 ;
        RECT 0 17.023 1.246 28.977 ;
        RECT 0 17 1.2 29 ;
      LAYER MET2 ;
        RECT 0 17 65 29 ;
        RECT 0 3.5 65 15.5 ;
        RECT 57.3 3.5 58.3 29 ;
        RECT 52.7 3.5 53.7 29 ;
        RECT 48.1 3.5 49.1 29 ;
        RECT 43.5 3.5 44.5 29 ;
        RECT 38.9 3.5 39.9 29 ;
        RECT 34.3 3.5 35.3 29 ;
        RECT 29.7 3.5 30.7 29 ;
        RECT 25.1 3.5 26.1 29 ;
        RECT 20.5 3.5 21.5 29 ;
        RECT 15.9 3.5 16.9 29 ;
        RECT 11.3 3.5 12.3 29 ;
        RECT 6.7 3.5 7.7 29 ;
        RECT 0 78.5 65 89.5 ;
    END
  END VSSIO
  OBS
    LAYER MET1 SPACING 0.09 ;
      RECT 0 -20 65 110 ;
    LAYER MET2 SPACING 0.1 ;
      RECT 58.475 107.675 65 110 ;
      RECT 0 107.675 6.525 110 ;
      RECT 0 107.675 65 108.825 ;
      RECT 0 -20 65 3.325 ;
      RECT 58.475 15.675 65 16.825 ;
      RECT 0 29.175 65 30.325 ;
      RECT 56.675 42.675 65 43.825 ;
      RECT 56.675 56.175 65 57.325 ;
      RECT 0 63.675 65 68.325 ;
      RECT 0 77.175 65 78.325 ;
      RECT 0 89.675 65 90.825 ;
      RECT 0 98.175 65 99.325 ;
      RECT 53.875 15.675 57.125 16.825 ;
      RECT 52.075 42.675 54.325 43.825 ;
      RECT 52.075 56.175 54.325 57.325 ;
      RECT 49.275 15.675 52.525 16.825 ;
      RECT 47.475 42.675 49.725 43.825 ;
      RECT 47.475 56.175 49.725 57.325 ;
      RECT 44.675 15.675 47.925 16.825 ;
      RECT 42.875 42.675 45.125 43.825 ;
      RECT 42.875 56.175 45.125 57.325 ;
      RECT 40.075 15.675 43.325 16.825 ;
      RECT 38.275 42.675 40.525 43.825 ;
      RECT 38.275 56.175 40.525 57.325 ;
      RECT 35.475 15.675 38.725 16.825 ;
      RECT 33.675 42.675 35.925 43.825 ;
      RECT 33.675 56.175 35.925 57.325 ;
      RECT 30.875 15.675 34.125 16.825 ;
      RECT 29.075 42.675 31.325 43.825 ;
      RECT 29.075 56.175 31.325 57.325 ;
      RECT 26.275 15.675 29.525 16.825 ;
      RECT 24.475 42.675 26.725 43.825 ;
      RECT 24.475 56.175 26.725 57.325 ;
      RECT 21.675 15.675 24.925 16.825 ;
      RECT 19.875 42.675 22.125 43.825 ;
      RECT 19.875 56.175 22.125 57.325 ;
      RECT 17.075 15.675 20.325 16.825 ;
      RECT 15.275 42.675 17.525 43.825 ;
      RECT 15.275 56.175 17.525 57.325 ;
      RECT 12.475 15.675 15.725 16.825 ;
      RECT 10.675 42.675 12.925 43.825 ;
      RECT 10.675 56.175 12.925 57.325 ;
      RECT 7.875 15.675 11.125 16.825 ;
      RECT 0 42.675 8.325 43.825 ;
      RECT 0 56.175 8.325 57.325 ;
      RECT 0 15.675 6.525 16.825 ;
    LAYER MET3 SPACING 0.1 ;
      RECT 0 63.675 65 68.325 ;
      RECT 1.375 63.665 65 68.325 ;
      RECT 3 57.5 62 68.325 ;
      RECT 57 -20 62 68.325 ;
      RECT 43 -20 50.5 68.325 ;
      RECT 29 -20 36.5 68.325 ;
      RECT 15 -20 22.5 68.325 ;
      RECT 3 -20 8.5 68.325 ;
      RECT 56.665 56.165 65 57.335 ;
      RECT 42.865 56.165 50.5 57.335 ;
      RECT 1.375 56.165 8.5 57.335 ;
      RECT 0 56.175 8.5 57.325 ;
      RECT 3 43.5 62 51 ;
      RECT 56.665 42.665 65 43.835 ;
      RECT 0 42.675 8.5 43.825 ;
      RECT 52.065 42.665 54.335 51 ;
      RECT 42.865 42.665 50.5 51 ;
      RECT 38.265 42.665 40.535 51 ;
      RECT 24.465 42.665 26.735 51 ;
      RECT 10.665 42.665 12.935 51 ;
      RECT 1.375 42.665 8.5 43.835 ;
      RECT 3 29.165 62 37 ;
      RECT 1.375 29.165 65 30.335 ;
      RECT 0 29.175 65 30.325 ;
      RECT 3 15.5 62 23 ;
      RECT 1.375 15.665 65 16.835 ;
      RECT 0 15.675 65 16.825 ;
      RECT 3 -20 62 9 ;
      RECT 1.375 -20 65 3.335 ;
      RECT 0 -20 65 3.325 ;
      RECT 63.8 3.5 65 15.5 ;
      RECT 63.776 3.512 65 15.488 ;
      RECT 63.73 3.547 65 15.453 ;
      RECT 63.684 3.593 65 15.407 ;
      RECT 63.638 3.639 65 15.361 ;
      RECT 63.592 3.685 65 15.315 ;
      RECT 63.546 3.731 65 15.269 ;
      RECT 63.5 3.777 65 15.223 ;
      RECT 63.8 17 65 29 ;
      RECT 63.776 17.012 65 28.988 ;
      RECT 63.73 17.047 65 28.953 ;
      RECT 63.684 17.093 65 28.907 ;
      RECT 63.638 17.139 65 28.861 ;
      RECT 63.592 17.185 65 28.815 ;
      RECT 63.546 17.231 65 28.769 ;
      RECT 63.5 17.277 65 28.723 ;
      RECT 63.8 30.5 65 42.5 ;
      RECT 63.776 30.512 65 42.488 ;
      RECT 63.73 30.547 65 42.453 ;
      RECT 63.684 30.593 65 42.407 ;
      RECT 63.638 30.639 65 42.361 ;
      RECT 63.592 30.685 65 42.315 ;
      RECT 63.546 30.731 65 42.269 ;
      RECT 63.5 30.777 65 42.223 ;
      RECT 63.8 44 65 56 ;
      RECT 63.776 44.012 65 55.988 ;
      RECT 63.73 44.047 65 55.953 ;
      RECT 63.684 44.093 65 55.907 ;
      RECT 63.638 44.139 65 55.861 ;
      RECT 63.592 44.185 65 55.815 ;
      RECT 63.546 44.231 65 55.769 ;
      RECT 63.5 44.277 65 55.723 ;
      RECT 63.8 57.5 65 63.5 ;
      RECT 63.776 57.512 65 63.488 ;
      RECT 63.73 57.547 65 63.453 ;
      RECT 63.684 57.593 65 63.407 ;
      RECT 63.638 57.639 65 63.361 ;
      RECT 63.592 57.685 65 63.315 ;
      RECT 63.546 57.731 65 63.269 ;
      RECT 63.5 57.777 65 63.223 ;
      RECT 58.475 107.675 65 110 ;
      RECT 0 107.675 6.525 110 ;
      RECT 0 107.675 65 108.825 ;
      RECT 0 77.175 65 78.325 ;
      RECT 0 89.675 65 90.825 ;
      RECT 0 98.175 65 99.325 ;
      RECT 52.065 56.165 54.335 57.335 ;
      RECT 38.265 56.165 40.535 57.335 ;
      RECT 24.465 56.165 26.735 57.335 ;
      RECT 10.665 56.165 12.935 57.335 ;
    LAYER MET4 SPACING 0.1 ;
      RECT 0 63.675 65 68.325 ;
      RECT 1.675 -20 65 68.325 ;
      RECT 1.375 63.652 65 68.325 ;
      RECT 1.651 63.387 65 68.325 ;
      RECT 1.421 63.606 65 68.325 ;
      RECT 1.605 63.422 65 68.325 ;
      RECT 1.467 63.56 65 68.325 ;
      RECT 1.559 63.468 65 68.325 ;
      RECT 1.513 63.514 65 68.325 ;
      RECT 1.651 55.887 65 57.613 ;
      RECT 1.605 55.922 65 57.578 ;
      RECT 1.559 55.968 65 57.532 ;
      RECT 1.513 56.014 65 57.486 ;
      RECT 1.467 56.06 65 57.44 ;
      RECT 1.421 56.106 65 57.394 ;
      RECT 1.375 56.152 65 57.348 ;
      RECT 0 56.175 65 57.325 ;
      RECT 1.651 42.387 65 44.113 ;
      RECT 1.605 42.422 65 44.078 ;
      RECT 1.559 42.468 65 44.032 ;
      RECT 1.513 42.514 65 43.986 ;
      RECT 1.467 42.56 65 43.94 ;
      RECT 1.421 42.606 65 43.894 ;
      RECT 1.375 42.652 65 43.848 ;
      RECT 0 42.675 65 43.825 ;
      RECT 1.651 28.887 65 30.613 ;
      RECT 1.605 28.922 65 30.578 ;
      RECT 1.559 28.968 65 30.532 ;
      RECT 1.513 29.014 65 30.486 ;
      RECT 1.467 29.06 65 30.44 ;
      RECT 1.421 29.106 65 30.394 ;
      RECT 1.375 29.152 65 30.348 ;
      RECT 0 29.175 65 30.325 ;
      RECT 1.651 15.387 65 17.113 ;
      RECT 1.605 15.422 65 17.078 ;
      RECT 1.559 15.468 65 17.032 ;
      RECT 1.513 15.514 65 16.986 ;
      RECT 1.467 15.56 65 16.94 ;
      RECT 1.421 15.606 65 16.894 ;
      RECT 1.375 15.652 65 16.848 ;
      RECT 0 15.675 65 16.825 ;
      RECT 1.651 -20 65 3.613 ;
      RECT 1.605 -20 65 3.578 ;
      RECT 1.559 -20 65 3.532 ;
      RECT 1.513 -20 65 3.486 ;
      RECT 1.467 -20 65 3.44 ;
      RECT 1.421 -20 65 3.394 ;
      RECT 1.375 -20 65 3.348 ;
      RECT 0 -20 65 3.325 ;
      RECT 58.475 107.675 65 110 ;
      RECT 0 107.675 6.525 110 ;
      RECT 0 107.675 65 108.825 ;
      RECT 0 77.175 65 78.325 ;
      RECT 0 89.675 65 90.825 ;
      RECT 0 98.175 65 99.325 ;
    LAYER MET5 SPACING 0.1 ;
      RECT 0 63.83 65 68.17 ;
      RECT 1.83 -20 65 68.17 ;
      RECT 1.53 63.807 65 68.17 ;
      RECT 1.806 63.542 65 68.17 ;
      RECT 1.576 63.761 65 68.17 ;
      RECT 1.76 63.577 65 68.17 ;
      RECT 1.622 63.715 65 68.17 ;
      RECT 1.714 63.623 65 68.17 ;
      RECT 1.668 63.669 65 68.17 ;
      RECT 1.806 56.042 65 57.458 ;
      RECT 1.76 56.077 65 57.423 ;
      RECT 1.714 56.123 65 57.377 ;
      RECT 1.668 56.169 65 57.331 ;
      RECT 1.622 56.215 65 57.285 ;
      RECT 1.576 56.261 65 57.239 ;
      RECT 1.53 56.307 65 57.193 ;
      RECT 0 56.33 65 57.17 ;
      RECT 1.806 42.542 65 43.958 ;
      RECT 1.76 42.577 65 43.923 ;
      RECT 1.714 42.623 65 43.877 ;
      RECT 1.668 42.669 65 43.831 ;
      RECT 1.622 42.715 65 43.785 ;
      RECT 1.576 42.761 65 43.739 ;
      RECT 1.53 42.807 65 43.693 ;
      RECT 0 42.83 65 43.67 ;
      RECT 1.806 29.042 65 30.458 ;
      RECT 1.76 29.077 65 30.423 ;
      RECT 1.714 29.123 65 30.377 ;
      RECT 1.668 29.169 65 30.331 ;
      RECT 1.622 29.215 65 30.285 ;
      RECT 1.576 29.261 65 30.239 ;
      RECT 1.53 29.307 65 30.193 ;
      RECT 0 29.33 65 30.17 ;
      RECT 1.806 15.542 65 16.958 ;
      RECT 1.76 15.577 65 16.923 ;
      RECT 1.714 15.623 65 16.877 ;
      RECT 1.668 15.669 65 16.831 ;
      RECT 1.622 15.715 65 16.785 ;
      RECT 1.576 15.761 65 16.739 ;
      RECT 1.53 15.807 65 16.693 ;
      RECT 0 15.83 65 16.67 ;
      RECT 1.806 -20 65 3.458 ;
      RECT 1.76 -20 65 3.423 ;
      RECT 1.714 -20 65 3.377 ;
      RECT 1.668 -20 65 3.331 ;
      RECT 1.622 -20 65 3.285 ;
      RECT 1.576 -20 65 3.239 ;
      RECT 1.53 -20 65 3.193 ;
      RECT 0 -20 65 3.17 ;
      RECT 58.63 107.83 65 110 ;
      RECT 0 107.83 6.37 110 ;
      RECT 0 107.83 65 108.67 ;
      RECT 0 77.33 65 78.17 ;
      RECT 0 89.83 65 90.67 ;
      RECT 0 98.33 65 99.17 ;
    LAYER T4M2 SPACING 0.4 ;
      RECT 64.584 -20 65 -3.193 ;
      RECT 0 -20 0.428 -3.205 ;
      RECT 64.538 -20 65 -3.239 ;
      RECT 0 -20 0.474 -3.251 ;
      RECT 64.492 -20 65 -3.285 ;
      RECT 0 -20 0.52 -3.297 ;
      RECT 64.446 -20 65 -3.331 ;
      RECT 0 -20 0.566 -3.343 ;
      RECT 64.4 -20 65 -3.377 ;
      RECT 0 -20 0.6 -3.383 ;
      RECT 0 -20 65 -3.4 ;
      RECT 58.9 108.1 65 110 ;
      RECT 0 108.1 6.1 110 ;
    LAYER RDL SPACING 2 ;
      RECT 0 -20 65 -5 ;
      RECT 0 72 65 110 ;
      RECT 3 4.5 62 63.5 ;
  END
END P65_1233_VSS1

MACRO P65_1233_VSS1A
  CLASS PAD ;
  ORIGIN 0 20 ;
  FOREIGN P65_1233_VSS1A 0 -20 ;
  SIZE 65 BY 130 ;
  SYMMETRY X Y R90 ;
  SITE IOSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET2 ;
        RECT 0 99.98 6.5 107.02 ;
        RECT 0 99.937 6.46 107.063 ;
        RECT 0 99.891 6.414 107.109 ;
        RECT 0 99.845 6.368 107.155 ;
        RECT 0 99.799 6.322 107.201 ;
        RECT 0 99.753 6.276 107.247 ;
        RECT 0 99.707 6.23 107.293 ;
        RECT 0 99.661 6.184 107.339 ;
        RECT 0 99.615 6.138 107.385 ;
        RECT 0 99.569 6.092 107.431 ;
        RECT 0 99.523 6.046 107.477 ;
        RECT 0 99.5 6 107.5 ;
    END
    PORT
      CLASS CORE ;
      LAYER MET5 ;
        RECT 0 99.5 65 107.5 ;
      LAYER MET4 ;
        RECT 0 99.5 65 107.5 ;
      LAYER MET3 ;
        RECT 0 99.5 65 107.5 ;
    END
  END VDD
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET5 ;
        RECT 0 68.5 65 77 ;
        RECT 0 30.788 1.5 42.212 ;
        RECT 0 30.753 1.476 42.247 ;
        RECT 0 30.707 1.43 42.293 ;
        RECT 0 30.661 1.384 42.339 ;
        RECT 0 30.615 1.338 42.385 ;
        RECT 0 30.569 1.292 42.431 ;
        RECT 0 30.523 1.246 42.477 ;
        RECT 0 30.5 1.2 42.5 ;
        RECT 0 44.288 1.5 55.712 ;
        RECT 0 44.253 1.476 55.747 ;
        RECT 0 44.207 1.43 55.793 ;
        RECT 0 44.161 1.384 55.839 ;
        RECT 0 44.115 1.338 55.885 ;
        RECT 0 44.069 1.292 55.931 ;
        RECT 0 44.023 1.246 55.977 ;
        RECT 0 44 1.2 56 ;
        RECT 0 57.788 1.5 63.212 ;
        RECT 0 57.753 1.476 63.247 ;
        RECT 0 57.707 1.43 63.293 ;
        RECT 0 57.661 1.384 63.339 ;
        RECT 0 57.615 1.338 63.385 ;
        RECT 0 57.569 1.292 63.431 ;
        RECT 0 57.523 1.246 63.477 ;
        RECT 0 57.5 1.2 63.5 ;
      LAYER MET4 ;
        RECT 0 68.5 65 77 ;
        RECT 0 30.788 1.5 42.212 ;
        RECT 0 30.753 1.476 42.247 ;
        RECT 0 30.707 1.43 42.293 ;
        RECT 0 30.661 1.384 42.339 ;
        RECT 0 30.615 1.338 42.385 ;
        RECT 0 30.569 1.292 42.431 ;
        RECT 0 30.523 1.246 42.477 ;
        RECT 0 30.5 1.2 42.5 ;
        RECT 0 44.288 1.5 55.712 ;
        RECT 0 44.253 1.476 55.747 ;
        RECT 0 44.207 1.43 55.793 ;
        RECT 0 44.161 1.384 55.839 ;
        RECT 0 44.115 1.338 55.885 ;
        RECT 0 44.069 1.292 55.931 ;
        RECT 0 44.023 1.246 55.977 ;
        RECT 0 44 1.2 56 ;
        RECT 0 57.788 1.5 63.212 ;
        RECT 0 57.753 1.476 63.247 ;
        RECT 0 57.707 1.43 63.293 ;
        RECT 0 57.661 1.384 63.339 ;
        RECT 0 57.615 1.338 63.385 ;
        RECT 0 57.569 1.292 63.431 ;
        RECT 0 57.523 1.246 63.477 ;
        RECT 0 57.5 1.2 63.5 ;
      LAYER MET3 ;
        RECT 0 68.5 65 77 ;
        RECT 0 30.788 1.5 42.212 ;
        RECT 0 30.753 1.476 42.247 ;
        RECT 0 30.707 1.43 42.293 ;
        RECT 0 30.661 1.384 42.339 ;
        RECT 0 30.615 1.338 42.385 ;
        RECT 0 30.569 1.292 42.431 ;
        RECT 0 30.523 1.246 42.477 ;
        RECT 0 30.5 1.2 42.5 ;
        RECT 0 44.288 1.5 55.712 ;
        RECT 0 44.253 1.476 55.747 ;
        RECT 0 44.207 1.43 55.793 ;
        RECT 0 44.161 1.384 55.839 ;
        RECT 0 44.115 1.338 55.885 ;
        RECT 0 44.069 1.292 55.931 ;
        RECT 0 44.023 1.246 55.977 ;
        RECT 0 44 1.2 56 ;
        RECT 0 57.788 1.5 63.212 ;
        RECT 0 57.753 1.476 63.247 ;
        RECT 0 57.707 1.43 63.293 ;
        RECT 0 57.661 1.384 63.339 ;
        RECT 0 57.615 1.338 63.385 ;
        RECT 0 57.569 1.292 63.431 ;
        RECT 0 57.523 1.246 63.477 ;
        RECT 0 57.5 1.2 63.5 ;
      LAYER MET2 ;
        RECT 0 57.5 65 63.5 ;
        RECT 0 44 65 56 ;
        RECT 0 30.5 65 42.5 ;
        RECT 56.015 30.5 59.205 63.5 ;
        RECT 50.435 30.5 53.625 63.5 ;
        RECT 44.855 30.5 48.045 63.5 ;
        RECT 39.275 30.5 42.465 63.5 ;
        RECT 33.695 30.5 36.885 63.5 ;
        RECT 28.115 30.5 31.305 63.5 ;
        RECT 22.535 30.5 25.725 63.5 ;
        RECT 16.955 30.5 20.145 63.5 ;
        RECT 11.375 30.5 14.565 63.5 ;
        RECT 5.795 30.5 8.985 63.5 ;
        RECT 0 68.98 6.5 76.52 ;
        RECT 0 68.937 6.46 76.563 ;
        RECT 0 68.891 6.414 76.609 ;
        RECT 0 68.845 6.368 76.655 ;
        RECT 0 68.799 6.322 76.701 ;
        RECT 0 68.753 6.276 76.747 ;
        RECT 0 68.707 6.23 76.793 ;
        RECT 0 68.661 6.184 76.839 ;
        RECT 0 68.615 6.138 76.885 ;
        RECT 0 68.569 6.092 76.931 ;
        RECT 0 68.523 6.046 76.977 ;
        RECT 0 68.5 6 77 ;
    END
  END VDDA
  PIN VSS
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 6.2694 LAYER VIA4 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 2.3085 LAYER VIA2 ;
    PORT
      LAYER MET5 ;
        RECT 0 91 65 98 ;
      LAYER MET4 ;
        RECT 0 91 65 98 ;
      LAYER MET3 ;
        RECT 0 91 65 98 ;
      LAYER MET2 ;
        RECT 0 91.48 6.5 97.52 ;
        RECT 0 91.437 6.46 97.563 ;
        RECT 0 91.391 6.414 97.609 ;
        RECT 0 91.345 6.368 97.655 ;
        RECT 0 91.299 6.322 97.701 ;
        RECT 0 91.253 6.276 97.747 ;
        RECT 0 91.207 6.23 97.793 ;
        RECT 0 91.161 6.184 97.839 ;
        RECT 0 91.115 6.138 97.885 ;
        RECT 0 91.069 6.092 97.931 ;
        RECT 0 91.023 6.046 97.977 ;
        RECT 0 91 6 98 ;
    END
  END VSS
  PIN VSSA
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA2 ;
    ANTENNAPARTIALCUTAREA 9.7524 LAYER VIA4 ;
    ANTENNAPARTIALCUTAREA 34.2144 LAYER T4V2 ;
    PORT
      LAYER T4M2 ;
        RECT 57 17 65 29 ;
        RECT 57 3.5 65 15.5 ;
        RECT 57 0.983 62 66.017 ;
        RECT 57 0.943 61.966 66.057 ;
        RECT 57 0.897 61.92 66.103 ;
        RECT 57 0.851 61.874 66.149 ;
        RECT 57 0.805 61.828 66.195 ;
        RECT 57 0.759 61.782 66.241 ;
        RECT 57 0.713 61.736 66.287 ;
        RECT 57 0.667 61.69 66.333 ;
        RECT 57 0.621 61.644 66.379 ;
        RECT 57 0.575 61.598 66.425 ;
        RECT 57 0.529 61.552 66.471 ;
        RECT 57 0.483 61.506 66.517 ;
        RECT 57 0.437 61.46 66.563 ;
        RECT 57 0.391 61.414 66.609 ;
        RECT 57 0.345 61.368 66.655 ;
        RECT 57 0.299 61.322 66.701 ;
        RECT 57 0.253 61.276 66.747 ;
        RECT 57 0.207 61.23 66.793 ;
        RECT 57 0.161 61.184 66.839 ;
        RECT 57 0.115 61.138 66.885 ;
        RECT 57 0.069 61.092 66.931 ;
        RECT 57 0.023 61.046 66.977 ;
        RECT 4 57.5 61 67 ;
        RECT 3 43.5 62 51 ;
        RECT 3 29.5 62 37 ;
        RECT 3 15.5 62 23 ;
        RECT 4 0 61 9 ;
        RECT 43 0 50.5 67 ;
        RECT 29 0 36.5 67 ;
        RECT 15 0 22.5 67 ;
        RECT 3 0.977 8.5 66.023 ;
        RECT 3.966 0.017 8.5 66.983 ;
        RECT 3.92 0.057 8.5 66.943 ;
        RECT 3.874 0.103 8.5 66.897 ;
        RECT 3.828 0.149 8.5 66.851 ;
        RECT 3.782 0.195 8.5 66.805 ;
        RECT 3.736 0.241 8.5 66.759 ;
        RECT 3.69 0.287 8.5 66.713 ;
        RECT 3.644 0.333 8.5 66.667 ;
        RECT 3.598 0.379 8.5 66.621 ;
        RECT 3.552 0.425 8.5 66.575 ;
        RECT 3.506 0.471 8.5 66.529 ;
        RECT 3.46 0.517 8.5 66.483 ;
        RECT 3.414 0.563 8.5 66.437 ;
        RECT 3.368 0.609 8.5 66.391 ;
        RECT 3.322 0.655 8.5 66.345 ;
        RECT 3.276 0.701 8.5 66.299 ;
        RECT 3.23 0.747 8.5 66.253 ;
        RECT 3.184 0.793 8.5 66.207 ;
        RECT 3.138 0.839 8.5 66.161 ;
        RECT 3.092 0.885 8.5 66.115 ;
        RECT 3.046 0.931 8.5 66.069 ;
        RECT 0 17 8.5 29 ;
        RECT 0 3.5 8.5 15.5 ;
      LAYER MET5 ;
        RECT 57 17 65 29 ;
        RECT 57 3.5 65 15.5 ;
        RECT 57 0.983 62 66.017 ;
        RECT 57 0.943 61.966 66.057 ;
        RECT 57 0.897 61.92 66.103 ;
        RECT 57 0.851 61.874 66.149 ;
        RECT 57 0.805 61.828 66.195 ;
        RECT 57 0.759 61.782 66.241 ;
        RECT 57 0.713 61.736 66.287 ;
        RECT 57 0.667 61.69 66.333 ;
        RECT 57 0.621 61.644 66.379 ;
        RECT 57 0.575 61.598 66.425 ;
        RECT 57 0.529 61.552 66.471 ;
        RECT 57 0.483 61.506 66.517 ;
        RECT 57 0.437 61.46 66.563 ;
        RECT 57 0.391 61.414 66.609 ;
        RECT 57 0.345 61.368 66.655 ;
        RECT 57 0.299 61.322 66.701 ;
        RECT 57 0.253 61.276 66.747 ;
        RECT 57 0.207 61.23 66.793 ;
        RECT 57 0.161 61.184 66.839 ;
        RECT 57 0.115 61.138 66.885 ;
        RECT 57 0.069 61.092 66.931 ;
        RECT 57 0.023 61.046 66.977 ;
        RECT 4 57.5 61 67 ;
        RECT 3 43.5 62 51 ;
        RECT 3 29.5 62 37 ;
        RECT 3 15.5 62 23 ;
        RECT 4 0 61 9 ;
        RECT 43 0 50.5 67 ;
        RECT 29 0 36.5 67 ;
        RECT 15 0 22.5 67 ;
        RECT 3 0.977 8.5 66.023 ;
        RECT 3.966 0.017 8.5 66.983 ;
        RECT 3.92 0.057 8.5 66.943 ;
        RECT 3.874 0.103 8.5 66.897 ;
        RECT 3.828 0.149 8.5 66.851 ;
        RECT 3.782 0.195 8.5 66.805 ;
        RECT 3.736 0.241 8.5 66.759 ;
        RECT 3.69 0.287 8.5 66.713 ;
        RECT 3.644 0.333 8.5 66.667 ;
        RECT 3.598 0.379 8.5 66.621 ;
        RECT 3.552 0.425 8.5 66.575 ;
        RECT 3.506 0.471 8.5 66.529 ;
        RECT 3.46 0.517 8.5 66.483 ;
        RECT 3.414 0.563 8.5 66.437 ;
        RECT 3.368 0.609 8.5 66.391 ;
        RECT 3.322 0.655 8.5 66.345 ;
        RECT 3.276 0.701 8.5 66.299 ;
        RECT 3.23 0.747 8.5 66.253 ;
        RECT 3.184 0.793 8.5 66.207 ;
        RECT 3.138 0.839 8.5 66.161 ;
        RECT 3.092 0.885 8.5 66.115 ;
        RECT 3.046 0.931 8.5 66.069 ;
        RECT 0 17 8.5 29 ;
        RECT 0 3.5 8.5 15.5 ;
        RECT 0 78.5 65 89.5 ;
        RECT 8 109 57 110 ;
      LAYER MET4 ;
        RECT 57 17 65 29 ;
        RECT 57 3.5 65 15.5 ;
        RECT 57 0.983 62 66.017 ;
        RECT 57 0.943 61.966 66.057 ;
        RECT 57 0.897 61.92 66.103 ;
        RECT 57 0.851 61.874 66.149 ;
        RECT 57 0.805 61.828 66.195 ;
        RECT 57 0.759 61.782 66.241 ;
        RECT 57 0.713 61.736 66.287 ;
        RECT 57 0.667 61.69 66.333 ;
        RECT 57 0.621 61.644 66.379 ;
        RECT 57 0.575 61.598 66.425 ;
        RECT 57 0.529 61.552 66.471 ;
        RECT 57 0.483 61.506 66.517 ;
        RECT 57 0.437 61.46 66.563 ;
        RECT 57 0.391 61.414 66.609 ;
        RECT 57 0.345 61.368 66.655 ;
        RECT 57 0.299 61.322 66.701 ;
        RECT 57 0.253 61.276 66.747 ;
        RECT 57 0.207 61.23 66.793 ;
        RECT 57 0.161 61.184 66.839 ;
        RECT 57 0.115 61.138 66.885 ;
        RECT 57 0.069 61.092 66.931 ;
        RECT 57 0.023 61.046 66.977 ;
        RECT 4 57.5 61 67 ;
        RECT 3 43.5 62 51 ;
        RECT 3 29.5 62 37 ;
        RECT 3 15.5 62 23 ;
        RECT 4 0 61 9 ;
        RECT 43 0 50.5 67 ;
        RECT 29 0 36.5 67 ;
        RECT 15 0 22.5 67 ;
        RECT 3 0.977 8.5 66.023 ;
        RECT 3.966 0.017 8.5 66.983 ;
        RECT 3.92 0.057 8.5 66.943 ;
        RECT 3.874 0.103 8.5 66.897 ;
        RECT 3.828 0.149 8.5 66.851 ;
        RECT 3.782 0.195 8.5 66.805 ;
        RECT 3.736 0.241 8.5 66.759 ;
        RECT 3.69 0.287 8.5 66.713 ;
        RECT 3.644 0.333 8.5 66.667 ;
        RECT 3.598 0.379 8.5 66.621 ;
        RECT 3.552 0.425 8.5 66.575 ;
        RECT 3.506 0.471 8.5 66.529 ;
        RECT 3.46 0.517 8.5 66.483 ;
        RECT 3.414 0.563 8.5 66.437 ;
        RECT 3.368 0.609 8.5 66.391 ;
        RECT 3.322 0.655 8.5 66.345 ;
        RECT 3.276 0.701 8.5 66.299 ;
        RECT 3.23 0.747 8.5 66.253 ;
        RECT 3.184 0.793 8.5 66.207 ;
        RECT 3.138 0.839 8.5 66.161 ;
        RECT 3.092 0.885 8.5 66.115 ;
        RECT 3.046 0.931 8.5 66.069 ;
        RECT 0 17 8.5 29 ;
        RECT 0 3.5 8.5 15.5 ;
        RECT 0 78.5 65 89.5 ;
        RECT 8 109 57 110 ;
      LAYER MET3 ;
        RECT 57 17 65 29 ;
        RECT 57 3.5 65 15.5 ;
        RECT 57 0.983 62 66.017 ;
        RECT 57 0.943 61.966 66.057 ;
        RECT 57 0.897 61.92 66.103 ;
        RECT 57 0.851 61.874 66.149 ;
        RECT 57 0.805 61.828 66.195 ;
        RECT 57 0.759 61.782 66.241 ;
        RECT 57 0.713 61.736 66.287 ;
        RECT 57 0.667 61.69 66.333 ;
        RECT 57 0.621 61.644 66.379 ;
        RECT 57 0.575 61.598 66.425 ;
        RECT 57 0.529 61.552 66.471 ;
        RECT 57 0.483 61.506 66.517 ;
        RECT 57 0.437 61.46 66.563 ;
        RECT 57 0.391 61.414 66.609 ;
        RECT 57 0.345 61.368 66.655 ;
        RECT 57 0.299 61.322 66.701 ;
        RECT 57 0.253 61.276 66.747 ;
        RECT 57 0.207 61.23 66.793 ;
        RECT 57 0.161 61.184 66.839 ;
        RECT 57 0.115 61.138 66.885 ;
        RECT 57 0.069 61.092 66.931 ;
        RECT 57 0.023 61.046 66.977 ;
        RECT 4 57.5 61 67 ;
        RECT 3 43.5 62 51 ;
        RECT 3 29.5 62 37 ;
        RECT 3 15.5 62 23 ;
        RECT 4 0 61 9 ;
        RECT 43 0 50.5 67 ;
        RECT 29 0 36.5 67 ;
        RECT 15 0 22.5 67 ;
        RECT 3 0.977 8.5 66.023 ;
        RECT 3.966 0.017 8.5 66.983 ;
        RECT 3.92 0.057 8.5 66.943 ;
        RECT 3.874 0.103 8.5 66.897 ;
        RECT 3.828 0.149 8.5 66.851 ;
        RECT 3.782 0.195 8.5 66.805 ;
        RECT 3.736 0.241 8.5 66.759 ;
        RECT 3.69 0.287 8.5 66.713 ;
        RECT 3.644 0.333 8.5 66.667 ;
        RECT 3.598 0.379 8.5 66.621 ;
        RECT 3.552 0.425 8.5 66.575 ;
        RECT 3.506 0.471 8.5 66.529 ;
        RECT 3.46 0.517 8.5 66.483 ;
        RECT 3.414 0.563 8.5 66.437 ;
        RECT 3.368 0.609 8.5 66.391 ;
        RECT 3.322 0.655 8.5 66.345 ;
        RECT 3.276 0.701 8.5 66.299 ;
        RECT 3.23 0.747 8.5 66.253 ;
        RECT 3.184 0.793 8.5 66.207 ;
        RECT 3.138 0.839 8.5 66.161 ;
        RECT 3.092 0.885 8.5 66.115 ;
        RECT 3.046 0.931 8.5 66.069 ;
        RECT 0 17 8.5 29 ;
        RECT 0 3.5 8.5 15.5 ;
        RECT 0 78.5 65 89.5 ;
        RECT 8 109 57 110 ;
      LAYER MET2 ;
        RECT 0 17 65 29 ;
        RECT 0 3.5 65 15.5 ;
        RECT 59.805 3.5 60.995 29 ;
        RECT 54.225 3.5 55.415 29 ;
        RECT 48.645 3.5 49.835 29 ;
        RECT 43.065 3.5 44.255 29 ;
        RECT 37.485 3.5 38.675 29 ;
        RECT 31.905 3.5 33.095 29 ;
        RECT 26.325 3.5 27.515 29 ;
        RECT 20.745 3.5 21.935 29 ;
        RECT 15.165 3.5 16.355 29 ;
        RECT 9.585 3.5 10.775 29 ;
        RECT 4.005 3.5 5.195 29 ;
        RECT 0 78.5 65 89.5 ;
        RECT 3 65 62 67 ;
        RECT 8 109 57 110 ;
        RECT 45.98 65 57 110 ;
        RECT 8 65 57 69.28 ;
        RECT 33.32 65 44.32 110 ;
        RECT 20.66 65 31.66 110 ;
        RECT 8 65 19 110 ;
    END
  END VSSA
  OBS
    LAYER MET1 SPACING 0.09 ;
      RECT 0 -20 65 110 ;
    LAYER MET2 SPACING 0.1 ;
      RECT 57.175 67.175 65 78.325 ;
      RECT 62.175 63.675 65 78.325 ;
      RECT 0 77.175 7.825 78.325 ;
      RECT 6.675 67.175 7.825 78.325 ;
      RECT 6.175 77.152 7.825 78.325 ;
      RECT 6.635 76.695 7.825 78.325 ;
      RECT 6.221 77.106 7.825 78.325 ;
      RECT 6.589 76.738 7.825 78.325 ;
      RECT 6.267 77.06 7.825 78.325 ;
      RECT 6.543 76.784 7.825 78.325 ;
      RECT 6.313 77.014 7.825 78.325 ;
      RECT 6.497 76.83 7.825 78.325 ;
      RECT 6.359 76.968 7.825 78.325 ;
      RECT 6.451 76.876 7.825 78.325 ;
      RECT 6.405 76.922 7.825 78.325 ;
      RECT 6.635 67.175 7.825 68.805 ;
      RECT 6.589 67.175 7.825 68.762 ;
      RECT 6.543 67.175 7.825 68.716 ;
      RECT 6.497 67.175 7.825 68.67 ;
      RECT 6.451 67.175 7.825 68.624 ;
      RECT 6.405 67.175 7.825 68.578 ;
      RECT 6.359 67.175 7.825 68.532 ;
      RECT 6.313 67.175 7.825 68.486 ;
      RECT 6.267 67.175 7.825 68.44 ;
      RECT 6.221 67.175 7.825 68.394 ;
      RECT 6.175 67.175 7.825 68.348 ;
      RECT 0 67.175 7.825 68.325 ;
      RECT 0 63.675 2.825 68.325 ;
      RECT 0 63.675 65 64.825 ;
      RECT 0 107.675 7.825 110 ;
      RECT 6.675 89.675 7.825 110 ;
      RECT 6.175 107.652 7.825 110 ;
      RECT 6.635 107.195 7.825 110 ;
      RECT 6.221 107.606 7.825 110 ;
      RECT 6.589 107.238 7.825 110 ;
      RECT 6.267 107.56 7.825 110 ;
      RECT 6.543 107.284 7.825 110 ;
      RECT 6.313 107.514 7.825 110 ;
      RECT 6.497 107.33 7.825 110 ;
      RECT 6.359 107.468 7.825 110 ;
      RECT 6.451 107.376 7.825 110 ;
      RECT 6.405 107.422 7.825 110 ;
      RECT 6.635 97.695 7.825 99.805 ;
      RECT 6.589 97.738 7.825 99.762 ;
      RECT 6.543 97.784 7.825 99.716 ;
      RECT 6.497 97.83 7.825 99.67 ;
      RECT 6.451 97.876 7.825 99.624 ;
      RECT 6.405 97.922 7.825 99.578 ;
      RECT 6.359 97.968 7.825 99.532 ;
      RECT 6.313 98.014 7.825 99.486 ;
      RECT 6.267 98.06 7.825 99.44 ;
      RECT 6.221 98.106 7.825 99.394 ;
      RECT 6.175 98.152 7.825 99.348 ;
      RECT 0 98.175 7.825 99.325 ;
      RECT 6.635 89.675 7.825 91.305 ;
      RECT 6.589 89.675 7.825 91.262 ;
      RECT 6.543 89.675 7.825 91.216 ;
      RECT 6.497 89.675 7.825 91.17 ;
      RECT 6.451 89.675 7.825 91.124 ;
      RECT 6.405 89.675 7.825 91.078 ;
      RECT 6.359 89.675 7.825 91.032 ;
      RECT 6.313 89.675 7.825 90.986 ;
      RECT 6.267 89.675 7.825 90.94 ;
      RECT 6.221 89.675 7.825 90.894 ;
      RECT 6.175 89.675 7.825 90.848 ;
      RECT 0 89.675 7.825 90.825 ;
      RECT 0 -20 65 3.325 ;
      RECT 61.17 15.675 65 16.825 ;
      RECT 0 29.175 65 30.325 ;
      RECT 59.38 42.675 65 43.825 ;
      RECT 59.38 56.175 65 57.325 ;
      RECT 57.175 89.675 65 110 ;
      RECT 55.59 15.675 59.63 16.825 ;
      RECT 53.8 42.675 55.84 43.825 ;
      RECT 53.8 56.175 55.84 57.325 ;
      RECT 50.01 15.675 54.05 16.825 ;
      RECT 48.22 42.675 50.26 43.825 ;
      RECT 48.22 56.175 50.26 57.325 ;
      RECT 44.43 15.675 48.47 16.825 ;
      RECT 44.495 69.455 45.805 78.325 ;
      RECT 44.495 89.675 45.805 108.825 ;
      RECT 42.64 42.675 44.68 43.825 ;
      RECT 42.64 56.175 44.68 57.325 ;
      RECT 38.85 15.675 42.89 16.825 ;
      RECT 37.06 42.675 39.1 43.825 ;
      RECT 37.06 56.175 39.1 57.325 ;
      RECT 33.27 15.675 37.31 16.825 ;
      RECT 31.48 42.675 33.52 43.825 ;
      RECT 31.48 56.175 33.52 57.325 ;
      RECT 31.835 69.455 33.145 78.325 ;
      RECT 31.835 89.675 33.145 108.825 ;
      RECT 27.69 15.675 31.73 16.825 ;
      RECT 25.9 42.675 27.94 43.825 ;
      RECT 25.9 56.175 27.94 57.325 ;
      RECT 22.11 15.675 26.15 16.825 ;
      RECT 20.32 42.675 22.36 43.825 ;
      RECT 20.32 56.175 22.36 57.325 ;
      RECT 16.53 15.675 20.57 16.825 ;
      RECT 19.175 69.455 20.485 78.325 ;
      RECT 19.175 89.675 20.485 108.825 ;
      RECT 14.74 42.675 16.78 43.825 ;
      RECT 14.74 56.175 16.78 57.325 ;
      RECT 10.95 15.675 14.99 16.825 ;
      RECT 9.16 42.675 11.2 43.825 ;
      RECT 9.16 56.175 11.2 57.325 ;
      RECT 5.37 15.675 9.41 16.825 ;
      RECT 0 42.675 5.62 43.825 ;
      RECT 0 56.175 5.62 57.325 ;
      RECT 0 15.675 3.83 16.825 ;
    LAYER MET3 SPACING 0.1 ;
      RECT 62.175 -20 65 3.325 ;
      RECT 0 -20 2.825 3.325 ;
      RECT 62.141 -20 65 0.808 ;
      RECT 0 -20 2.871 0.802 ;
      RECT 62.095 -20 65 0.768 ;
      RECT 0 -20 2.917 0.756 ;
      RECT 62.049 -20 65 0.722 ;
      RECT 0 -20 2.963 0.71 ;
      RECT 62.003 -20 65 0.676 ;
      RECT 0 -20 3.009 0.664 ;
      RECT 61.957 -20 65 0.63 ;
      RECT 0 -20 3.055 0.618 ;
      RECT 61.911 -20 65 0.584 ;
      RECT 0 -20 3.101 0.572 ;
      RECT 61.865 -20 65 0.538 ;
      RECT 0 -20 3.147 0.526 ;
      RECT 61.819 -20 65 0.492 ;
      RECT 0 -20 3.193 0.48 ;
      RECT 61.773 -20 65 0.446 ;
      RECT 0 -20 3.239 0.434 ;
      RECT 61.727 -20 65 0.4 ;
      RECT 0 -20 3.285 0.388 ;
      RECT 61.681 -20 65 0.354 ;
      RECT 0 -20 3.331 0.342 ;
      RECT 61.635 -20 65 0.308 ;
      RECT 0 -20 3.377 0.296 ;
      RECT 61.589 -20 65 0.262 ;
      RECT 0 -20 3.423 0.25 ;
      RECT 61.543 -20 65 0.216 ;
      RECT 0 -20 3.469 0.204 ;
      RECT 61.497 -20 65 0.17 ;
      RECT 0 -20 3.515 0.158 ;
      RECT 61.451 -20 65 0.124 ;
      RECT 0 -20 3.561 0.112 ;
      RECT 61.405 -20 65 0.078 ;
      RECT 0 -20 3.607 0.066 ;
      RECT 61.359 -20 65 0.032 ;
      RECT 0 -20 3.653 0.02 ;
      RECT 61.313 -20 65 -0.014 ;
      RECT 0 -20 3.699 -0.026 ;
      RECT 61.267 -20 65 -0.06 ;
      RECT 0 -20 3.745 -0.072 ;
      RECT 61.221 -20 65 -0.106 ;
      RECT 0 -20 3.791 -0.118 ;
      RECT 61.175 -20 65 -0.152 ;
      RECT 0 -20 3.825 -0.158 ;
      RECT 0 -20 65 -0.175 ;
      RECT 63.8 30.5 65 42.5 ;
      RECT 63.776 30.512 65 42.488 ;
      RECT 63.73 30.547 65 42.453 ;
      RECT 63.684 30.593 65 42.407 ;
      RECT 63.638 30.639 65 42.361 ;
      RECT 63.592 30.685 65 42.315 ;
      RECT 63.546 30.731 65 42.269 ;
      RECT 63.5 30.777 65 42.223 ;
      RECT 63.8 44 65 56 ;
      RECT 63.776 44.012 65 55.988 ;
      RECT 63.73 44.047 65 55.953 ;
      RECT 63.684 44.093 65 55.907 ;
      RECT 63.638 44.139 65 55.861 ;
      RECT 63.592 44.185 65 55.815 ;
      RECT 63.546 44.231 65 55.769 ;
      RECT 63.5 44.277 65 55.723 ;
      RECT 63.8 57.5 65 63.5 ;
      RECT 63.776 57.512 65 63.488 ;
      RECT 63.73 57.547 65 63.453 ;
      RECT 63.684 57.593 65 63.407 ;
      RECT 63.638 57.639 65 63.361 ;
      RECT 63.592 57.685 65 63.315 ;
      RECT 63.546 57.731 65 63.269 ;
      RECT 63.5 57.777 65 63.223 ;
      RECT 57.165 67.175 65 68.325 ;
      RECT 62.175 63.665 65 68.325 ;
      RECT 61.175 67.165 65 68.325 ;
      RECT 62.165 66.192 65 68.325 ;
      RECT 57.175 107.675 65 110 ;
      RECT 57.165 107.675 65 108.825 ;
      RECT 0 67.175 7.835 68.325 ;
      RECT 0 67.165 3.825 68.325 ;
      RECT 0 66.198 2.835 68.325 ;
      RECT 0 63.675 2.825 68.325 ;
      RECT 1.375 63.665 2.825 68.325 ;
      RECT 0 107.675 7.825 110 ;
      RECT 0 107.675 7.835 108.825 ;
      RECT 1.375 29.175 2.825 30.335 ;
      RECT 0 29.175 2.825 30.325 ;
      RECT 1.375 42.665 2.825 43.835 ;
      RECT 0 42.675 2.825 43.825 ;
      RECT 1.375 56.165 2.825 57.335 ;
      RECT 0 56.175 2.825 57.325 ;
      RECT 62.175 15.675 65 16.825 ;
      RECT 62.175 29.175 65 30.335 ;
      RECT 62.175 42.665 65 43.835 ;
      RECT 62.175 56.165 65 57.335 ;
      RECT 57.165 77.175 65 78.325 ;
      RECT 57.165 89.675 65 90.825 ;
      RECT 57.165 98.175 65 99.325 ;
      RECT 50.675 29.165 56.825 29.325 ;
      RECT 53.79 42.665 55.85 43.325 ;
      RECT 53.79 56.165 55.85 57.325 ;
      RECT 44.485 77.175 45.815 78.325 ;
      RECT 44.485 89.675 45.815 90.825 ;
      RECT 44.485 98.175 45.815 99.325 ;
      RECT 44.485 107.675 45.815 108.825 ;
      RECT 36.675 29.165 42.825 29.325 ;
      RECT 42.63 42.665 42.825 43.325 ;
      RECT 42.63 56.165 42.825 57.325 ;
      RECT 37.05 42.665 39.11 43.325 ;
      RECT 37.05 56.165 39.11 57.325 ;
      RECT 31.825 77.175 33.155 78.325 ;
      RECT 31.825 89.675 33.155 90.825 ;
      RECT 31.825 98.175 33.155 99.325 ;
      RECT 31.825 107.675 33.155 108.825 ;
      RECT 22.675 29.165 28.825 29.325 ;
      RECT 25.89 42.665 27.95 43.325 ;
      RECT 25.89 56.165 27.95 57.325 ;
      RECT 19.165 77.175 20.495 78.325 ;
      RECT 19.165 89.675 20.495 90.825 ;
      RECT 19.165 98.175 20.495 99.325 ;
      RECT 19.165 107.675 20.495 108.825 ;
      RECT 8.675 29.165 14.825 29.325 ;
      RECT 9.15 42.665 11.21 43.325 ;
      RECT 9.15 56.165 11.21 57.325 ;
      RECT 0 77.175 7.835 78.325 ;
      RECT 0 89.675 7.835 90.825 ;
      RECT 0 98.175 7.835 99.325 ;
      RECT 0 15.675 2.825 16.825 ;
    LAYER MET4 SPACING 0.1 ;
      RECT 62.175 -20 65 3.325 ;
      RECT 0 -20 2.825 3.325 ;
      RECT 62.141 -20 65 0.808 ;
      RECT 0 -20 2.871 0.802 ;
      RECT 62.095 -20 65 0.768 ;
      RECT 0 -20 2.917 0.756 ;
      RECT 62.049 -20 65 0.722 ;
      RECT 0 -20 2.963 0.71 ;
      RECT 62.003 -20 65 0.676 ;
      RECT 0 -20 3.009 0.664 ;
      RECT 61.957 -20 65 0.63 ;
      RECT 0 -20 3.055 0.618 ;
      RECT 61.911 -20 65 0.584 ;
      RECT 0 -20 3.101 0.572 ;
      RECT 61.865 -20 65 0.538 ;
      RECT 0 -20 3.147 0.526 ;
      RECT 61.819 -20 65 0.492 ;
      RECT 0 -20 3.193 0.48 ;
      RECT 61.773 -20 65 0.446 ;
      RECT 0 -20 3.239 0.434 ;
      RECT 61.727 -20 65 0.4 ;
      RECT 0 -20 3.285 0.388 ;
      RECT 61.681 -20 65 0.354 ;
      RECT 0 -20 3.331 0.342 ;
      RECT 61.635 -20 65 0.308 ;
      RECT 0 -20 3.377 0.296 ;
      RECT 61.589 -20 65 0.262 ;
      RECT 0 -20 3.423 0.25 ;
      RECT 61.543 -20 65 0.216 ;
      RECT 0 -20 3.469 0.204 ;
      RECT 61.497 -20 65 0.17 ;
      RECT 0 -20 3.515 0.158 ;
      RECT 61.451 -20 65 0.124 ;
      RECT 0 -20 3.561 0.112 ;
      RECT 61.405 -20 65 0.078 ;
      RECT 0 -20 3.607 0.066 ;
      RECT 61.359 -20 65 0.032 ;
      RECT 0 -20 3.653 0.02 ;
      RECT 61.313 -20 65 -0.014 ;
      RECT 0 -20 3.699 -0.026 ;
      RECT 61.267 -20 65 -0.06 ;
      RECT 0 -20 3.745 -0.072 ;
      RECT 61.221 -20 65 -0.106 ;
      RECT 0 -20 3.791 -0.118 ;
      RECT 61.175 -20 65 -0.152 ;
      RECT 0 -20 3.825 -0.158 ;
      RECT 0 -20 65 -0.175 ;
      RECT 0 67.175 65 68.325 ;
      RECT 62.175 29.175 65 68.325 ;
      RECT 61.175 67.152 65 68.325 ;
      RECT 62.141 66.192 65 68.325 ;
      RECT 0 67.158 3.825 68.325 ;
      RECT 0 67.118 3.791 68.325 ;
      RECT 61.221 67.106 65 68.325 ;
      RECT 62.095 66.232 65 68.325 ;
      RECT 0 67.072 3.745 68.325 ;
      RECT 61.267 67.06 65 68.325 ;
      RECT 62.049 66.278 65 68.325 ;
      RECT 0 67.026 3.699 68.325 ;
      RECT 61.313 67.014 65 68.325 ;
      RECT 62.003 66.324 65 68.325 ;
      RECT 0 66.98 3.653 68.325 ;
      RECT 61.359 66.968 65 68.325 ;
      RECT 61.957 66.37 65 68.325 ;
      RECT 0 66.934 3.607 68.325 ;
      RECT 61.405 66.922 65 68.325 ;
      RECT 61.911 66.416 65 68.325 ;
      RECT 0 66.888 3.561 68.325 ;
      RECT 61.451 66.876 65 68.325 ;
      RECT 61.865 66.462 65 68.325 ;
      RECT 0 66.842 3.515 68.325 ;
      RECT 61.497 66.83 65 68.325 ;
      RECT 61.819 66.508 65 68.325 ;
      RECT 0 66.796 3.469 68.325 ;
      RECT 61.543 66.784 65 68.325 ;
      RECT 61.773 66.554 65 68.325 ;
      RECT 0 66.75 3.423 68.325 ;
      RECT 61.589 66.738 65 68.325 ;
      RECT 61.727 66.6 65 68.325 ;
      RECT 0 66.704 3.377 68.325 ;
      RECT 61.635 66.692 65 68.325 ;
      RECT 61.681 66.646 65 68.325 ;
      RECT 0 66.658 3.331 68.325 ;
      RECT 0 66.612 3.285 68.325 ;
      RECT 0 66.566 3.239 68.325 ;
      RECT 0 66.52 3.193 68.325 ;
      RECT 0 66.474 3.147 68.325 ;
      RECT 0 66.428 3.101 68.325 ;
      RECT 0 66.382 3.055 68.325 ;
      RECT 0 66.336 3.009 68.325 ;
      RECT 0 66.29 2.963 68.325 ;
      RECT 0 66.244 2.917 68.325 ;
      RECT 0 66.198 2.871 68.325 ;
      RECT 0 63.675 2.825 68.325 ;
      RECT 1.675 29.175 2.825 68.325 ;
      RECT 1.375 63.652 2.825 68.325 ;
      RECT 1.651 63.387 2.825 68.325 ;
      RECT 1.421 63.606 2.825 68.325 ;
      RECT 1.605 63.422 2.825 68.325 ;
      RECT 1.467 63.56 2.825 68.325 ;
      RECT 1.559 63.468 2.825 68.325 ;
      RECT 1.513 63.514 2.825 68.325 ;
      RECT 1.651 55.887 2.825 57.613 ;
      RECT 1.605 55.922 2.825 57.578 ;
      RECT 1.559 55.968 2.825 57.532 ;
      RECT 1.513 56.014 2.825 57.486 ;
      RECT 1.467 56.06 2.825 57.44 ;
      RECT 1.421 56.106 2.825 57.394 ;
      RECT 1.375 56.152 2.825 57.348 ;
      RECT 0 56.175 2.825 57.325 ;
      RECT 1.651 42.387 2.825 44.113 ;
      RECT 1.605 42.422 2.825 44.078 ;
      RECT 1.559 42.468 2.825 44.032 ;
      RECT 1.513 42.514 2.825 43.986 ;
      RECT 1.467 42.56 2.825 43.94 ;
      RECT 1.421 42.606 2.825 43.894 ;
      RECT 1.375 42.652 2.825 43.848 ;
      RECT 0 42.675 2.825 43.825 ;
      RECT 1.651 29.175 2.825 30.613 ;
      RECT 1.605 29.175 2.825 30.578 ;
      RECT 1.559 29.175 2.825 30.532 ;
      RECT 1.513 29.175 2.825 30.486 ;
      RECT 1.467 29.175 2.825 30.44 ;
      RECT 1.421 29.175 2.825 30.394 ;
      RECT 1.375 29.175 2.825 30.348 ;
      RECT 0 29.175 2.825 30.325 ;
      RECT 57.175 107.675 65 110 ;
      RECT 0 107.675 7.825 110 ;
      RECT 0 107.675 65 108.825 ;
      RECT 62.175 15.675 65 16.825 ;
      RECT 0 77.175 65 78.325 ;
      RECT 0 89.675 65 90.825 ;
      RECT 0 98.175 65 99.325 ;
      RECT 50.675 9.175 56.825 15.325 ;
      RECT 50.675 23.175 56.825 29.325 ;
      RECT 50.675 37.175 56.825 43.325 ;
      RECT 50.675 51.175 56.825 57.325 ;
      RECT 36.675 9.175 42.825 15.325 ;
      RECT 36.675 23.175 42.825 29.325 ;
      RECT 36.675 37.175 42.825 43.325 ;
      RECT 36.675 51.175 42.825 57.325 ;
      RECT 22.675 9.175 28.825 15.325 ;
      RECT 22.675 23.175 28.825 29.325 ;
      RECT 22.675 37.175 28.825 43.325 ;
      RECT 22.675 51.175 28.825 57.325 ;
      RECT 8.675 9.175 14.825 15.325 ;
      RECT 8.675 23.175 14.825 29.325 ;
      RECT 8.675 37.175 14.825 43.325 ;
      RECT 8.675 51.175 14.825 57.325 ;
      RECT 0 15.675 2.825 16.825 ;
    LAYER MET5 SPACING 0.1 ;
      RECT 62.33 -20 65 3.17 ;
      RECT 0 -20 2.67 3.17 ;
      RECT 62.296 -20 65 0.653 ;
      RECT 0 -20 2.716 0.647 ;
      RECT 62.25 -20 65 0.613 ;
      RECT 0 -20 2.762 0.601 ;
      RECT 62.204 -20 65 0.567 ;
      RECT 0 -20 2.808 0.555 ;
      RECT 62.158 -20 65 0.521 ;
      RECT 0 -20 2.854 0.509 ;
      RECT 62.112 -20 65 0.475 ;
      RECT 0 -20 2.9 0.463 ;
      RECT 62.066 -20 65 0.429 ;
      RECT 0 -20 2.946 0.417 ;
      RECT 62.02 -20 65 0.383 ;
      RECT 0 -20 2.992 0.371 ;
      RECT 61.974 -20 65 0.337 ;
      RECT 0 -20 3.038 0.325 ;
      RECT 61.928 -20 65 0.291 ;
      RECT 0 -20 3.084 0.279 ;
      RECT 61.882 -20 65 0.245 ;
      RECT 0 -20 3.13 0.233 ;
      RECT 61.836 -20 65 0.199 ;
      RECT 0 -20 3.176 0.187 ;
      RECT 61.79 -20 65 0.153 ;
      RECT 0 -20 3.222 0.141 ;
      RECT 61.744 -20 65 0.107 ;
      RECT 0 -20 3.268 0.095 ;
      RECT 61.698 -20 65 0.061 ;
      RECT 0 -20 3.314 0.049 ;
      RECT 61.652 -20 65 0.015 ;
      RECT 0 -20 3.36 0.003 ;
      RECT 61.606 -20 65 -0.031 ;
      RECT 0 -20 3.406 -0.043 ;
      RECT 61.56 -20 65 -0.077 ;
      RECT 0 -20 3.452 -0.089 ;
      RECT 61.514 -20 65 -0.123 ;
      RECT 0 -20 3.498 -0.135 ;
      RECT 61.468 -20 65 -0.169 ;
      RECT 0 -20 3.544 -0.181 ;
      RECT 61.422 -20 65 -0.215 ;
      RECT 0 -20 3.59 -0.227 ;
      RECT 61.376 -20 65 -0.261 ;
      RECT 0 -20 3.636 -0.273 ;
      RECT 61.33 -20 65 -0.307 ;
      RECT 0 -20 3.67 -0.313 ;
      RECT 0 -20 65 -0.33 ;
      RECT 0 67.33 65 68.17 ;
      RECT 62.33 29.33 65 68.17 ;
      RECT 61.33 67.307 65 68.17 ;
      RECT 62.296 66.347 65 68.17 ;
      RECT 0 67.313 3.67 68.17 ;
      RECT 0 67.273 3.636 68.17 ;
      RECT 61.376 67.261 65 68.17 ;
      RECT 62.25 66.387 65 68.17 ;
      RECT 0 67.227 3.59 68.17 ;
      RECT 61.422 67.215 65 68.17 ;
      RECT 62.204 66.433 65 68.17 ;
      RECT 0 67.181 3.544 68.17 ;
      RECT 61.468 67.169 65 68.17 ;
      RECT 62.158 66.479 65 68.17 ;
      RECT 0 67.135 3.498 68.17 ;
      RECT 61.514 67.123 65 68.17 ;
      RECT 62.112 66.525 65 68.17 ;
      RECT 0 67.089 3.452 68.17 ;
      RECT 61.56 67.077 65 68.17 ;
      RECT 62.066 66.571 65 68.17 ;
      RECT 0 67.043 3.406 68.17 ;
      RECT 61.606 67.031 65 68.17 ;
      RECT 62.02 66.617 65 68.17 ;
      RECT 0 66.997 3.36 68.17 ;
      RECT 61.652 66.985 65 68.17 ;
      RECT 61.974 66.663 65 68.17 ;
      RECT 0 66.951 3.314 68.17 ;
      RECT 61.698 66.939 65 68.17 ;
      RECT 61.928 66.709 65 68.17 ;
      RECT 0 66.905 3.268 68.17 ;
      RECT 61.744 66.893 65 68.17 ;
      RECT 61.882 66.755 65 68.17 ;
      RECT 0 66.859 3.222 68.17 ;
      RECT 61.79 66.847 65 68.17 ;
      RECT 61.836 66.801 65 68.17 ;
      RECT 0 66.813 3.176 68.17 ;
      RECT 0 66.767 3.13 68.17 ;
      RECT 0 66.721 3.084 68.17 ;
      RECT 0 66.675 3.038 68.17 ;
      RECT 0 66.629 2.992 68.17 ;
      RECT 0 66.583 2.946 68.17 ;
      RECT 0 66.537 2.9 68.17 ;
      RECT 0 66.491 2.854 68.17 ;
      RECT 0 66.445 2.808 68.17 ;
      RECT 0 66.399 2.762 68.17 ;
      RECT 0 66.353 2.716 68.17 ;
      RECT 0 63.83 2.67 68.17 ;
      RECT 1.83 29.33 2.67 68.17 ;
      RECT 1.53 63.807 2.67 68.17 ;
      RECT 1.806 63.542 2.67 68.17 ;
      RECT 1.576 63.761 2.67 68.17 ;
      RECT 1.76 63.577 2.67 68.17 ;
      RECT 1.622 63.715 2.67 68.17 ;
      RECT 1.714 63.623 2.67 68.17 ;
      RECT 1.668 63.669 2.67 68.17 ;
      RECT 1.806 56.042 2.67 57.458 ;
      RECT 1.76 56.077 2.67 57.423 ;
      RECT 1.714 56.123 2.67 57.377 ;
      RECT 1.668 56.169 2.67 57.331 ;
      RECT 1.622 56.215 2.67 57.285 ;
      RECT 1.576 56.261 2.67 57.239 ;
      RECT 1.53 56.307 2.67 57.193 ;
      RECT 0 56.33 2.67 57.17 ;
      RECT 1.806 42.542 2.67 43.958 ;
      RECT 1.76 42.577 2.67 43.923 ;
      RECT 1.714 42.623 2.67 43.877 ;
      RECT 1.668 42.669 2.67 43.831 ;
      RECT 1.622 42.715 2.67 43.785 ;
      RECT 1.576 42.761 2.67 43.739 ;
      RECT 1.53 42.807 2.67 43.693 ;
      RECT 0 42.83 2.67 43.67 ;
      RECT 1.806 29.33 2.67 30.458 ;
      RECT 1.76 29.33 2.67 30.423 ;
      RECT 1.714 29.33 2.67 30.377 ;
      RECT 1.668 29.33 2.67 30.331 ;
      RECT 1.622 29.33 2.67 30.285 ;
      RECT 1.576 29.33 2.67 30.239 ;
      RECT 1.53 29.33 2.67 30.193 ;
      RECT 0 29.33 2.67 30.17 ;
      RECT 57.33 107.83 65 110 ;
      RECT 0 107.83 7.67 110 ;
      RECT 0 107.83 65 108.67 ;
      RECT 62.33 15.83 65 16.67 ;
      RECT 0 77.33 65 78.17 ;
      RECT 0 89.83 65 90.67 ;
      RECT 0 98.33 65 99.17 ;
      RECT 50.83 9.33 56.67 15.17 ;
      RECT 50.83 23.33 56.67 29.17 ;
      RECT 50.83 37.33 56.67 43.17 ;
      RECT 50.83 51.33 56.67 57.17 ;
      RECT 36.83 9.33 42.67 15.17 ;
      RECT 36.83 23.33 42.67 29.17 ;
      RECT 36.83 37.33 42.67 43.17 ;
      RECT 36.83 51.33 42.67 57.17 ;
      RECT 22.83 9.33 28.67 15.17 ;
      RECT 22.83 23.33 28.67 29.17 ;
      RECT 22.83 37.33 28.67 43.17 ;
      RECT 22.83 51.33 28.67 57.17 ;
      RECT 8.83 9.33 14.67 15.17 ;
      RECT 8.83 23.33 14.67 29.17 ;
      RECT 8.83 37.33 14.67 43.17 ;
      RECT 8.83 51.33 14.67 57.17 ;
      RECT 0 15.83 2.67 16.67 ;
    LAYER T4M2 SPACING 0.4 ;
      RECT 64.584 -20 65 -3.193 ;
      RECT 0 -20 0.428 -3.205 ;
      RECT 64.538 -20 65 -3.239 ;
      RECT 0 -20 0.474 -3.251 ;
      RECT 64.492 -20 65 -3.285 ;
      RECT 0 -20 0.52 -3.297 ;
      RECT 64.446 -20 65 -3.331 ;
      RECT 0 -20 0.566 -3.343 ;
      RECT 64.4 -20 65 -3.377 ;
      RECT 0 -20 0.6 -3.383 ;
      RECT 0 -20 65 -3.4 ;
      RECT 57.6 108.1 65 110 ;
      RECT 0 108.1 7.4 110 ;
    LAYER RDL SPACING 2 ;
      RECT 0 -20 65 -5 ;
      RECT 0 72 65 110 ;
      RECT 3.5 5 61.5 63 ;
  END
END P65_1233_VSS1A

MACRO P65_1233_VSS3
  CLASS PAD ;
  ORIGIN 0 20 ;
  FOREIGN P65_1233_VSS3 0 -20 ;
  SIZE 65 BY 130 ;
  SYMMETRY X Y R90 ;
  SITE IOSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER MET5 ;
        RECT 0 99.5 65 107.5 ;
      LAYER MET4 ;
        RECT 0 99.5 65 107.5 ;
      LAYER MET3 ;
        RECT 0 99.5 65 107.5 ;
      LAYER MET2 ;
        RECT 0 99.5 65 107.5 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET5 ;
        RECT 0 68.5 65 77 ;
        RECT 0 30.788 1.5 42.212 ;
        RECT 0 30.753 1.476 42.247 ;
        RECT 0 30.707 1.43 42.293 ;
        RECT 0 30.661 1.384 42.339 ;
        RECT 0 30.615 1.338 42.385 ;
        RECT 0 30.569 1.292 42.431 ;
        RECT 0 30.523 1.246 42.477 ;
        RECT 0 30.5 1.2 42.5 ;
        RECT 0 44.288 1.5 55.712 ;
        RECT 0 44.253 1.476 55.747 ;
        RECT 0 44.207 1.43 55.793 ;
        RECT 0 44.161 1.384 55.839 ;
        RECT 0 44.115 1.338 55.885 ;
        RECT 0 44.069 1.292 55.931 ;
        RECT 0 44.023 1.246 55.977 ;
        RECT 0 44 1.2 56 ;
        RECT 0 57.788 1.5 63.212 ;
        RECT 0 57.753 1.476 63.247 ;
        RECT 0 57.707 1.43 63.293 ;
        RECT 0 57.661 1.384 63.339 ;
        RECT 0 57.615 1.338 63.385 ;
        RECT 0 57.569 1.292 63.431 ;
        RECT 0 57.523 1.246 63.477 ;
        RECT 0 57.5 1.2 63.5 ;
      LAYER MET4 ;
        RECT 0 68.5 65 77 ;
        RECT 0 30.788 1.5 42.212 ;
        RECT 0 30.753 1.476 42.247 ;
        RECT 0 30.707 1.43 42.293 ;
        RECT 0 30.661 1.384 42.339 ;
        RECT 0 30.615 1.338 42.385 ;
        RECT 0 30.569 1.292 42.431 ;
        RECT 0 30.523 1.246 42.477 ;
        RECT 0 30.5 1.2 42.5 ;
        RECT 0 44.288 1.5 55.712 ;
        RECT 0 44.253 1.476 55.747 ;
        RECT 0 44.207 1.43 55.793 ;
        RECT 0 44.161 1.384 55.839 ;
        RECT 0 44.115 1.338 55.885 ;
        RECT 0 44.069 1.292 55.931 ;
        RECT 0 44.023 1.246 55.977 ;
        RECT 0 44 1.2 56 ;
        RECT 0 57.788 1.5 63.212 ;
        RECT 0 57.753 1.476 63.247 ;
        RECT 0 57.707 1.43 63.293 ;
        RECT 0 57.661 1.384 63.339 ;
        RECT 0 57.615 1.338 63.385 ;
        RECT 0 57.569 1.292 63.431 ;
        RECT 0 57.523 1.246 63.477 ;
        RECT 0 57.5 1.2 63.5 ;
      LAYER MET3 ;
        RECT 0 68.5 65 77 ;
        RECT 0 30.788 1.5 42.212 ;
        RECT 0 30.753 1.476 42.247 ;
        RECT 0 30.707 1.43 42.293 ;
        RECT 0 30.661 1.384 42.339 ;
        RECT 0 30.615 1.338 42.385 ;
        RECT 0 30.569 1.292 42.431 ;
        RECT 0 30.523 1.246 42.477 ;
        RECT 0 30.5 1.2 42.5 ;
        RECT 0 44.288 1.5 55.712 ;
        RECT 0 44.253 1.476 55.747 ;
        RECT 0 44.207 1.43 55.793 ;
        RECT 0 44.161 1.384 55.839 ;
        RECT 0 44.115 1.338 55.885 ;
        RECT 0 44.069 1.292 55.931 ;
        RECT 0 44.023 1.246 55.977 ;
        RECT 0 44 1.2 56 ;
        RECT 0 57.788 1.5 63.212 ;
        RECT 0 57.753 1.476 63.247 ;
        RECT 0 57.707 1.43 63.293 ;
        RECT 0 57.661 1.384 63.339 ;
        RECT 0 57.615 1.338 63.385 ;
        RECT 0 57.569 1.292 63.431 ;
        RECT 0 57.523 1.246 63.477 ;
        RECT 0 57.5 1.2 63.5 ;
      LAYER MET2 ;
        RECT 0 57.5 65 63.5 ;
        RECT 0 44 65 56 ;
        RECT 0 30.5 65 42.5 ;
        RECT 54.5 30.5 56.5 63.5 ;
        RECT 49.9 30.5 51.9 63.5 ;
        RECT 45.3 30.5 47.3 63.5 ;
        RECT 40.7 30.5 42.7 63.5 ;
        RECT 36.1 30.5 38.1 63.5 ;
        RECT 31.5 30.5 33.5 63.5 ;
        RECT 26.9 30.5 28.9 63.5 ;
        RECT 22.3 30.5 24.3 63.5 ;
        RECT 17.7 30.5 19.7 63.5 ;
        RECT 13.1 30.5 15.1 63.5 ;
        RECT 8.5 30.5 10.5 63.5 ;
        RECT 0 68.5 65 77 ;
    END
  END VDDIO
  PIN VSS
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3275 LAYER MET4 ;
    ANTENNAPARTIALMETALAREA 3275 LAYER MET3 ;
    ANTENNAPARTIALMETALAREA 3275 LAYER MET5 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 6.237 LAYER VIA2 ;
    ANTENNAPARTIALCUTAREA 6.2694 LAYER VIA4 ;
    ANTENNAPARTIALCUTAREA 34.992 LAYER T4V2 ;
    PORT
      LAYER T4M2 ;
        RECT 57 0.983 62 66.017 ;
        RECT 57 0.943 61.966 66.057 ;
        RECT 57 0.897 61.92 66.103 ;
        RECT 57 0.851 61.874 66.149 ;
        RECT 57 0.805 61.828 66.195 ;
        RECT 57 0.759 61.782 66.241 ;
        RECT 57 0.713 61.736 66.287 ;
        RECT 57 0.667 61.69 66.333 ;
        RECT 57 0.621 61.644 66.379 ;
        RECT 57 0.575 61.598 66.425 ;
        RECT 57 0.529 61.552 66.471 ;
        RECT 57 0.483 61.506 66.517 ;
        RECT 57 0.437 61.46 66.563 ;
        RECT 57 0.391 61.414 66.609 ;
        RECT 57 0.345 61.368 66.655 ;
        RECT 57 0.299 61.322 66.701 ;
        RECT 57 0.253 61.276 66.747 ;
        RECT 57 0.207 61.23 66.793 ;
        RECT 57 0.161 61.184 66.839 ;
        RECT 57 0.115 61.138 66.885 ;
        RECT 57 0.069 61.092 66.931 ;
        RECT 57 0.023 61.046 66.977 ;
        RECT 4 57.5 61 67 ;
        RECT 3 43.5 62 51 ;
        RECT 3 29.5 62 37 ;
        RECT 3 15.5 62 23 ;
        RECT 4 0 61 9 ;
        RECT 43 0 50.5 67 ;
        RECT 29 0 36.5 67 ;
        RECT 15 0 22.5 67 ;
        RECT 3 0.977 8.5 66.023 ;
        RECT 3.966 0.017 8.5 66.983 ;
        RECT 3.92 0.057 8.5 66.943 ;
        RECT 3.874 0.103 8.5 66.897 ;
        RECT 3.828 0.149 8.5 66.851 ;
        RECT 3.782 0.195 8.5 66.805 ;
        RECT 3.736 0.241 8.5 66.759 ;
        RECT 3.69 0.287 8.5 66.713 ;
        RECT 3.644 0.333 8.5 66.667 ;
        RECT 3.598 0.379 8.5 66.621 ;
        RECT 3.552 0.425 8.5 66.575 ;
        RECT 3.506 0.471 8.5 66.529 ;
        RECT 3.46 0.517 8.5 66.483 ;
        RECT 3.414 0.563 8.5 66.437 ;
        RECT 3.368 0.609 8.5 66.391 ;
        RECT 3.322 0.655 8.5 66.345 ;
        RECT 3.276 0.701 8.5 66.299 ;
        RECT 3.23 0.747 8.5 66.253 ;
        RECT 3.184 0.793 8.5 66.207 ;
        RECT 3.138 0.839 8.5 66.161 ;
        RECT 3.092 0.885 8.5 66.115 ;
        RECT 3.046 0.931 8.5 66.069 ;
      LAYER MET5 ;
        RECT 0 91 65 98 ;
        RECT 6.7 109 58.3 110 ;
      LAYER MET4 ;
        RECT 0 91 65 98 ;
        RECT 6.7 109 58.3 110 ;
      LAYER MET3 ;
        RECT 0 91 65 98 ;
        RECT 6.7 109 58.3 110 ;
      LAYER MET2 ;
        RECT 0 91 65 98 ;
        RECT 6.7 109 58.3 110 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA2 ;
    ANTENNAPARTIALCUTAREA 9.7524 LAYER VIA4 ;
    PORT
      LAYER MET5 ;
        RECT 0 78.5 65 89.5 ;
        RECT 0 3.788 1.5 15.212 ;
        RECT 0 3.753 1.476 15.247 ;
        RECT 0 3.707 1.43 15.293 ;
        RECT 0 3.661 1.384 15.339 ;
        RECT 0 3.615 1.338 15.385 ;
        RECT 0 3.569 1.292 15.431 ;
        RECT 0 3.523 1.246 15.477 ;
        RECT 0 3.5 1.2 15.5 ;
        RECT 0 17.288 1.5 28.712 ;
        RECT 0 17.253 1.476 28.747 ;
        RECT 0 17.207 1.43 28.793 ;
        RECT 0 17.161 1.384 28.839 ;
        RECT 0 17.115 1.338 28.885 ;
        RECT 0 17.069 1.292 28.931 ;
        RECT 0 17.023 1.246 28.977 ;
        RECT 0 17 1.2 29 ;
      LAYER MET4 ;
        RECT 0 78.5 65 89.5 ;
        RECT 0 3.788 1.5 15.212 ;
        RECT 0 3.753 1.476 15.247 ;
        RECT 0 3.707 1.43 15.293 ;
        RECT 0 3.661 1.384 15.339 ;
        RECT 0 3.615 1.338 15.385 ;
        RECT 0 3.569 1.292 15.431 ;
        RECT 0 3.523 1.246 15.477 ;
        RECT 0 3.5 1.2 15.5 ;
        RECT 0 17.288 1.5 28.712 ;
        RECT 0 17.253 1.476 28.747 ;
        RECT 0 17.207 1.43 28.793 ;
        RECT 0 17.161 1.384 28.839 ;
        RECT 0 17.115 1.338 28.885 ;
        RECT 0 17.069 1.292 28.931 ;
        RECT 0 17.023 1.246 28.977 ;
        RECT 0 17 1.2 29 ;
      LAYER MET3 ;
        RECT 0 78.5 65 89.5 ;
        RECT 0 3.788 1.5 15.212 ;
        RECT 0 3.753 1.476 15.247 ;
        RECT 0 3.707 1.43 15.293 ;
        RECT 0 3.661 1.384 15.339 ;
        RECT 0 3.615 1.338 15.385 ;
        RECT 0 3.569 1.292 15.431 ;
        RECT 0 3.523 1.246 15.477 ;
        RECT 0 3.5 1.2 15.5 ;
        RECT 0 17.288 1.5 28.712 ;
        RECT 0 17.253 1.476 28.747 ;
        RECT 0 17.207 1.43 28.793 ;
        RECT 0 17.161 1.384 28.839 ;
        RECT 0 17.115 1.338 28.885 ;
        RECT 0 17.069 1.292 28.931 ;
        RECT 0 17.023 1.246 28.977 ;
        RECT 0 17 1.2 29 ;
      LAYER MET2 ;
        RECT 0 17 65 29 ;
        RECT 0 3.5 65 15.5 ;
        RECT 57.3 3.5 58.3 29 ;
        RECT 52.7 3.5 53.7 29 ;
        RECT 48.1 3.5 49.1 29 ;
        RECT 43.5 3.5 44.5 29 ;
        RECT 38.9 3.5 39.9 29 ;
        RECT 34.3 3.5 35.3 29 ;
        RECT 29.7 3.5 30.7 29 ;
        RECT 25.1 3.5 26.1 29 ;
        RECT 20.5 3.5 21.5 29 ;
        RECT 15.9 3.5 16.9 29 ;
        RECT 11.3 3.5 12.3 29 ;
        RECT 6.7 3.5 7.7 29 ;
        RECT 0 78.5 65 89.5 ;
    END
  END VSSIO
  OBS
    LAYER MET1 SPACING 0.09 ;
      RECT 0 -20 65 110 ;
    LAYER MET2 SPACING 0.1 ;
      RECT 58.475 107.675 65 110 ;
      RECT 0 107.675 6.525 110 ;
      RECT 0 107.675 65 108.825 ;
      RECT 0 -20 65 3.325 ;
      RECT 58.475 15.675 65 16.825 ;
      RECT 0 29.175 65 30.325 ;
      RECT 56.675 42.675 65 43.825 ;
      RECT 56.675 56.175 65 57.325 ;
      RECT 0 63.675 65 68.325 ;
      RECT 0 77.175 65 78.325 ;
      RECT 0 89.675 65 90.825 ;
      RECT 0 98.175 65 99.325 ;
      RECT 53.875 15.675 57.125 16.825 ;
      RECT 52.075 42.675 54.325 43.825 ;
      RECT 52.075 56.175 54.325 57.325 ;
      RECT 49.275 15.675 52.525 16.825 ;
      RECT 47.475 42.675 49.725 43.825 ;
      RECT 47.475 56.175 49.725 57.325 ;
      RECT 44.675 15.675 47.925 16.825 ;
      RECT 42.875 42.675 45.125 43.825 ;
      RECT 42.875 56.175 45.125 57.325 ;
      RECT 40.075 15.675 43.325 16.825 ;
      RECT 38.275 42.675 40.525 43.825 ;
      RECT 38.275 56.175 40.525 57.325 ;
      RECT 35.475 15.675 38.725 16.825 ;
      RECT 33.675 42.675 35.925 43.825 ;
      RECT 33.675 56.175 35.925 57.325 ;
      RECT 30.875 15.675 34.125 16.825 ;
      RECT 29.075 42.675 31.325 43.825 ;
      RECT 29.075 56.175 31.325 57.325 ;
      RECT 26.275 15.675 29.525 16.825 ;
      RECT 24.475 42.675 26.725 43.825 ;
      RECT 24.475 56.175 26.725 57.325 ;
      RECT 21.675 15.675 24.925 16.825 ;
      RECT 19.875 42.675 22.125 43.825 ;
      RECT 19.875 56.175 22.125 57.325 ;
      RECT 17.075 15.675 20.325 16.825 ;
      RECT 15.275 42.675 17.525 43.825 ;
      RECT 15.275 56.175 17.525 57.325 ;
      RECT 12.475 15.675 15.725 16.825 ;
      RECT 10.675 42.675 12.925 43.825 ;
      RECT 10.675 56.175 12.925 57.325 ;
      RECT 7.875 15.675 11.125 16.825 ;
      RECT 0 42.675 8.325 43.825 ;
      RECT 0 56.175 8.325 57.325 ;
      RECT 0 15.675 6.525 16.825 ;
    LAYER MET3 SPACING 0.1 ;
      RECT 0 63.675 65 68.325 ;
      RECT 1.375 63.665 65 68.325 ;
      RECT 3 57.5 62 68.325 ;
      RECT 57 -20 62 68.325 ;
      RECT 43 -20 50.5 68.325 ;
      RECT 29 -20 36.5 68.325 ;
      RECT 15 -20 22.5 68.325 ;
      RECT 3 -20 8.5 68.325 ;
      RECT 56.665 56.165 65 57.335 ;
      RECT 42.865 56.165 50.5 57.335 ;
      RECT 1.375 56.165 8.5 57.335 ;
      RECT 0 56.175 8.5 57.325 ;
      RECT 3 43.5 62 51 ;
      RECT 56.665 42.665 65 43.835 ;
      RECT 0 42.675 8.5 43.825 ;
      RECT 52.065 42.665 54.335 51 ;
      RECT 42.865 42.665 50.5 51 ;
      RECT 38.265 42.665 40.535 51 ;
      RECT 24.465 42.665 26.735 51 ;
      RECT 10.665 42.665 12.935 51 ;
      RECT 1.375 42.665 8.5 43.835 ;
      RECT 3 29.165 62 37 ;
      RECT 1.375 29.165 65 30.335 ;
      RECT 0 29.175 65 30.325 ;
      RECT 3 15.5 62 23 ;
      RECT 1.375 15.665 65 16.835 ;
      RECT 0 15.675 65 16.825 ;
      RECT 3 -20 62 9 ;
      RECT 1.375 -20 65 3.335 ;
      RECT 0 -20 65 3.325 ;
      RECT 63.8 3.5 65 15.5 ;
      RECT 63.776 3.512 65 15.488 ;
      RECT 63.73 3.547 65 15.453 ;
      RECT 63.684 3.593 65 15.407 ;
      RECT 63.638 3.639 65 15.361 ;
      RECT 63.592 3.685 65 15.315 ;
      RECT 63.546 3.731 65 15.269 ;
      RECT 63.5 3.777 65 15.223 ;
      RECT 63.8 17 65 29 ;
      RECT 63.776 17.012 65 28.988 ;
      RECT 63.73 17.047 65 28.953 ;
      RECT 63.684 17.093 65 28.907 ;
      RECT 63.638 17.139 65 28.861 ;
      RECT 63.592 17.185 65 28.815 ;
      RECT 63.546 17.231 65 28.769 ;
      RECT 63.5 17.277 65 28.723 ;
      RECT 63.8 30.5 65 42.5 ;
      RECT 63.776 30.512 65 42.488 ;
      RECT 63.73 30.547 65 42.453 ;
      RECT 63.684 30.593 65 42.407 ;
      RECT 63.638 30.639 65 42.361 ;
      RECT 63.592 30.685 65 42.315 ;
      RECT 63.546 30.731 65 42.269 ;
      RECT 63.5 30.777 65 42.223 ;
      RECT 63.8 44 65 56 ;
      RECT 63.776 44.012 65 55.988 ;
      RECT 63.73 44.047 65 55.953 ;
      RECT 63.684 44.093 65 55.907 ;
      RECT 63.638 44.139 65 55.861 ;
      RECT 63.592 44.185 65 55.815 ;
      RECT 63.546 44.231 65 55.769 ;
      RECT 63.5 44.277 65 55.723 ;
      RECT 63.8 57.5 65 63.5 ;
      RECT 63.776 57.512 65 63.488 ;
      RECT 63.73 57.547 65 63.453 ;
      RECT 63.684 57.593 65 63.407 ;
      RECT 63.638 57.639 65 63.361 ;
      RECT 63.592 57.685 65 63.315 ;
      RECT 63.546 57.731 65 63.269 ;
      RECT 63.5 57.777 65 63.223 ;
      RECT 58.475 107.675 65 110 ;
      RECT 0 107.675 6.525 110 ;
      RECT 0 107.675 65 108.825 ;
      RECT 0 77.175 65 78.325 ;
      RECT 0 89.675 65 90.825 ;
      RECT 0 98.175 65 99.325 ;
      RECT 52.065 56.165 54.335 57.335 ;
      RECT 38.265 56.165 40.535 57.335 ;
      RECT 24.465 56.165 26.735 57.335 ;
      RECT 10.665 56.165 12.935 57.335 ;
    LAYER MET4 SPACING 0.1 ;
      RECT 0 63.675 65 68.325 ;
      RECT 1.675 -20 65 68.325 ;
      RECT 1.375 63.652 65 68.325 ;
      RECT 1.651 63.387 65 68.325 ;
      RECT 1.421 63.606 65 68.325 ;
      RECT 1.605 63.422 65 68.325 ;
      RECT 1.467 63.56 65 68.325 ;
      RECT 1.559 63.468 65 68.325 ;
      RECT 1.513 63.514 65 68.325 ;
      RECT 1.651 55.887 65 57.613 ;
      RECT 1.605 55.922 65 57.578 ;
      RECT 1.559 55.968 65 57.532 ;
      RECT 1.513 56.014 65 57.486 ;
      RECT 1.467 56.06 65 57.44 ;
      RECT 1.421 56.106 65 57.394 ;
      RECT 1.375 56.152 65 57.348 ;
      RECT 0 56.175 65 57.325 ;
      RECT 1.651 42.387 65 44.113 ;
      RECT 1.605 42.422 65 44.078 ;
      RECT 1.559 42.468 65 44.032 ;
      RECT 1.513 42.514 65 43.986 ;
      RECT 1.467 42.56 65 43.94 ;
      RECT 1.421 42.606 65 43.894 ;
      RECT 1.375 42.652 65 43.848 ;
      RECT 0 42.675 65 43.825 ;
      RECT 1.651 28.887 65 30.613 ;
      RECT 1.605 28.922 65 30.578 ;
      RECT 1.559 28.968 65 30.532 ;
      RECT 1.513 29.014 65 30.486 ;
      RECT 1.467 29.06 65 30.44 ;
      RECT 1.421 29.106 65 30.394 ;
      RECT 1.375 29.152 65 30.348 ;
      RECT 0 29.175 65 30.325 ;
      RECT 1.651 15.387 65 17.113 ;
      RECT 1.605 15.422 65 17.078 ;
      RECT 1.559 15.468 65 17.032 ;
      RECT 1.513 15.514 65 16.986 ;
      RECT 1.467 15.56 65 16.94 ;
      RECT 1.421 15.606 65 16.894 ;
      RECT 1.375 15.652 65 16.848 ;
      RECT 0 15.675 65 16.825 ;
      RECT 1.651 -20 65 3.613 ;
      RECT 1.605 -20 65 3.578 ;
      RECT 1.559 -20 65 3.532 ;
      RECT 1.513 -20 65 3.486 ;
      RECT 1.467 -20 65 3.44 ;
      RECT 1.421 -20 65 3.394 ;
      RECT 1.375 -20 65 3.348 ;
      RECT 0 -20 65 3.325 ;
      RECT 58.475 107.675 65 110 ;
      RECT 0 107.675 6.525 110 ;
      RECT 0 107.675 65 108.825 ;
      RECT 0 77.175 65 78.325 ;
      RECT 0 89.675 65 90.825 ;
      RECT 0 98.175 65 99.325 ;
    LAYER MET5 SPACING 0.1 ;
      RECT 0 63.83 65 68.17 ;
      RECT 1.83 -20 65 68.17 ;
      RECT 1.53 63.807 65 68.17 ;
      RECT 1.806 63.542 65 68.17 ;
      RECT 1.576 63.761 65 68.17 ;
      RECT 1.76 63.577 65 68.17 ;
      RECT 1.622 63.715 65 68.17 ;
      RECT 1.714 63.623 65 68.17 ;
      RECT 1.668 63.669 65 68.17 ;
      RECT 1.806 56.042 65 57.458 ;
      RECT 1.76 56.077 65 57.423 ;
      RECT 1.714 56.123 65 57.377 ;
      RECT 1.668 56.169 65 57.331 ;
      RECT 1.622 56.215 65 57.285 ;
      RECT 1.576 56.261 65 57.239 ;
      RECT 1.53 56.307 65 57.193 ;
      RECT 0 56.33 65 57.17 ;
      RECT 1.806 42.542 65 43.958 ;
      RECT 1.76 42.577 65 43.923 ;
      RECT 1.714 42.623 65 43.877 ;
      RECT 1.668 42.669 65 43.831 ;
      RECT 1.622 42.715 65 43.785 ;
      RECT 1.576 42.761 65 43.739 ;
      RECT 1.53 42.807 65 43.693 ;
      RECT 0 42.83 65 43.67 ;
      RECT 1.806 29.042 65 30.458 ;
      RECT 1.76 29.077 65 30.423 ;
      RECT 1.714 29.123 65 30.377 ;
      RECT 1.668 29.169 65 30.331 ;
      RECT 1.622 29.215 65 30.285 ;
      RECT 1.576 29.261 65 30.239 ;
      RECT 1.53 29.307 65 30.193 ;
      RECT 0 29.33 65 30.17 ;
      RECT 1.806 15.542 65 16.958 ;
      RECT 1.76 15.577 65 16.923 ;
      RECT 1.714 15.623 65 16.877 ;
      RECT 1.668 15.669 65 16.831 ;
      RECT 1.622 15.715 65 16.785 ;
      RECT 1.576 15.761 65 16.739 ;
      RECT 1.53 15.807 65 16.693 ;
      RECT 0 15.83 65 16.67 ;
      RECT 1.806 -20 65 3.458 ;
      RECT 1.76 -20 65 3.423 ;
      RECT 1.714 -20 65 3.377 ;
      RECT 1.668 -20 65 3.331 ;
      RECT 1.622 -20 65 3.285 ;
      RECT 1.576 -20 65 3.239 ;
      RECT 1.53 -20 65 3.193 ;
      RECT 0 -20 65 3.17 ;
      RECT 58.63 107.83 65 110 ;
      RECT 0 107.83 6.37 110 ;
      RECT 0 107.83 65 108.67 ;
      RECT 0 77.33 65 78.17 ;
      RECT 0 89.83 65 90.67 ;
      RECT 0 98.33 65 99.17 ;
    LAYER T4M2 SPACING 0.4 ;
      RECT 64.584 -20 65 -3.193 ;
      RECT 0 -20 0.428 -3.205 ;
      RECT 64.538 -20 65 -3.239 ;
      RECT 0 -20 0.474 -3.251 ;
      RECT 64.492 -20 65 -3.285 ;
      RECT 0 -20 0.52 -3.297 ;
      RECT 64.446 -20 65 -3.331 ;
      RECT 0 -20 0.566 -3.343 ;
      RECT 64.4 -20 65 -3.377 ;
      RECT 0 -20 0.6 -3.383 ;
      RECT 0 -20 65 -3.4 ;
      RECT 58.9 108.1 65 110 ;
      RECT 0 108.1 6.1 110 ;
    LAYER RDL SPACING 2 ;
      RECT 0 -20 65 -5 ;
      RECT 0 72 65 110 ;
      RECT 3 4.5 62 63.5 ;
  END
END P65_1233_VSS3

MACRO P65_1233_VSSIO3
  CLASS PAD ;
  ORIGIN 0 20 ;
  FOREIGN P65_1233_VSSIO3 0 -20 ;
  SIZE 65 BY 130 ;
  SYMMETRY X Y R90 ;
  SITE IOSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET2 ;
        RECT 0 99.98 6.5 107.02 ;
        RECT 0 99.937 6.46 107.063 ;
        RECT 0 99.891 6.414 107.109 ;
        RECT 0 99.845 6.368 107.155 ;
        RECT 0 99.799 6.322 107.201 ;
        RECT 0 99.753 6.276 107.247 ;
        RECT 0 99.707 6.23 107.293 ;
        RECT 0 99.661 6.184 107.339 ;
        RECT 0 99.615 6.138 107.385 ;
        RECT 0 99.569 6.092 107.431 ;
        RECT 0 99.523 6.046 107.477 ;
        RECT 0 99.5 6 107.5 ;
    END
    PORT
      CLASS CORE ;
      LAYER MET5 ;
        RECT 0 99.5 65 107.5 ;
      LAYER MET4 ;
        RECT 0 99.5 65 107.5 ;
      LAYER MET3 ;
        RECT 0 99.5 65 107.5 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET5 ;
        RECT 0 68.5 65 77 ;
        RECT 0 30.788 1.5 42.212 ;
        RECT 0 30.753 1.476 42.247 ;
        RECT 0 30.707 1.43 42.293 ;
        RECT 0 30.661 1.384 42.339 ;
        RECT 0 30.615 1.338 42.385 ;
        RECT 0 30.569 1.292 42.431 ;
        RECT 0 30.523 1.246 42.477 ;
        RECT 0 30.5 1.2 42.5 ;
        RECT 0 44.288 1.5 55.712 ;
        RECT 0 44.253 1.476 55.747 ;
        RECT 0 44.207 1.43 55.793 ;
        RECT 0 44.161 1.384 55.839 ;
        RECT 0 44.115 1.338 55.885 ;
        RECT 0 44.069 1.292 55.931 ;
        RECT 0 44.023 1.246 55.977 ;
        RECT 0 44 1.2 56 ;
        RECT 0 57.788 1.5 63.212 ;
        RECT 0 57.753 1.476 63.247 ;
        RECT 0 57.707 1.43 63.293 ;
        RECT 0 57.661 1.384 63.339 ;
        RECT 0 57.615 1.338 63.385 ;
        RECT 0 57.569 1.292 63.431 ;
        RECT 0 57.523 1.246 63.477 ;
        RECT 0 57.5 1.2 63.5 ;
      LAYER MET4 ;
        RECT 0 68.5 65 77 ;
        RECT 0 30.788 1.5 42.212 ;
        RECT 0 30.753 1.476 42.247 ;
        RECT 0 30.707 1.43 42.293 ;
        RECT 0 30.661 1.384 42.339 ;
        RECT 0 30.615 1.338 42.385 ;
        RECT 0 30.569 1.292 42.431 ;
        RECT 0 30.523 1.246 42.477 ;
        RECT 0 30.5 1.2 42.5 ;
        RECT 0 44.288 1.5 55.712 ;
        RECT 0 44.253 1.476 55.747 ;
        RECT 0 44.207 1.43 55.793 ;
        RECT 0 44.161 1.384 55.839 ;
        RECT 0 44.115 1.338 55.885 ;
        RECT 0 44.069 1.292 55.931 ;
        RECT 0 44.023 1.246 55.977 ;
        RECT 0 44 1.2 56 ;
        RECT 0 57.788 1.5 63.212 ;
        RECT 0 57.753 1.476 63.247 ;
        RECT 0 57.707 1.43 63.293 ;
        RECT 0 57.661 1.384 63.339 ;
        RECT 0 57.615 1.338 63.385 ;
        RECT 0 57.569 1.292 63.431 ;
        RECT 0 57.523 1.246 63.477 ;
        RECT 0 57.5 1.2 63.5 ;
      LAYER MET3 ;
        RECT 0 68.5 65 77 ;
        RECT 0 30.788 1.5 42.212 ;
        RECT 0 30.753 1.476 42.247 ;
        RECT 0 30.707 1.43 42.293 ;
        RECT 0 30.661 1.384 42.339 ;
        RECT 0 30.615 1.338 42.385 ;
        RECT 0 30.569 1.292 42.431 ;
        RECT 0 30.523 1.246 42.477 ;
        RECT 0 30.5 1.2 42.5 ;
        RECT 0 44.288 1.5 55.712 ;
        RECT 0 44.253 1.476 55.747 ;
        RECT 0 44.207 1.43 55.793 ;
        RECT 0 44.161 1.384 55.839 ;
        RECT 0 44.115 1.338 55.885 ;
        RECT 0 44.069 1.292 55.931 ;
        RECT 0 44.023 1.246 55.977 ;
        RECT 0 44 1.2 56 ;
        RECT 0 57.788 1.5 63.212 ;
        RECT 0 57.753 1.476 63.247 ;
        RECT 0 57.707 1.43 63.293 ;
        RECT 0 57.661 1.384 63.339 ;
        RECT 0 57.615 1.338 63.385 ;
        RECT 0 57.569 1.292 63.431 ;
        RECT 0 57.523 1.246 63.477 ;
        RECT 0 57.5 1.2 63.5 ;
      LAYER MET2 ;
        RECT 0 57.5 65 63.5 ;
        RECT 0 44 65 56 ;
        RECT 0 30.5 65 42.5 ;
        RECT 56.015 30.5 59.205 63.5 ;
        RECT 50.435 30.5 53.625 63.5 ;
        RECT 44.855 30.5 48.045 63.5 ;
        RECT 39.275 30.5 42.465 63.5 ;
        RECT 33.695 30.5 36.885 63.5 ;
        RECT 28.115 30.5 31.305 63.5 ;
        RECT 22.535 30.5 25.725 63.5 ;
        RECT 16.955 30.5 20.145 63.5 ;
        RECT 11.375 30.5 14.565 63.5 ;
        RECT 5.795 30.5 8.985 63.5 ;
        RECT 0 68.98 6.5 76.52 ;
        RECT 0 68.937 6.46 76.563 ;
        RECT 0 68.891 6.414 76.609 ;
        RECT 0 68.845 6.368 76.655 ;
        RECT 0 68.799 6.322 76.701 ;
        RECT 0 68.753 6.276 76.747 ;
        RECT 0 68.707 6.23 76.793 ;
        RECT 0 68.661 6.184 76.839 ;
        RECT 0 68.615 6.138 76.885 ;
        RECT 0 68.569 6.092 76.931 ;
        RECT 0 68.523 6.046 76.977 ;
        RECT 0 68.5 6 77 ;
    END
  END VDDIO
  PIN VSS
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 6.2694 LAYER VIA4 ;
    ANTENNAPARTIALCUTAREA 0.0081 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 2.3085 LAYER VIA2 ;
    PORT
      LAYER MET5 ;
        RECT 0 91 65 98 ;
      LAYER MET4 ;
        RECT 0 91 65 98 ;
      LAYER MET3 ;
        RECT 0 91 65 98 ;
      LAYER MET2 ;
        RECT 0 91.48 6.5 97.52 ;
        RECT 0 91.437 6.46 97.563 ;
        RECT 0 91.391 6.414 97.609 ;
        RECT 0 91.345 6.368 97.655 ;
        RECT 0 91.299 6.322 97.701 ;
        RECT 0 91.253 6.276 97.747 ;
        RECT 0 91.207 6.23 97.793 ;
        RECT 0 91.161 6.184 97.839 ;
        RECT 0 91.115 6.138 97.885 ;
        RECT 0 91.069 6.092 97.931 ;
        RECT 0 91.023 6.046 97.977 ;
        RECT 0 91 6 98 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 520 LAYER RDL ;
    ANTENNAPARTIALCUTAREA 5.85 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 5.85 LAYER VIA2 ;
    ANTENNAPARTIALCUTAREA 9.7524 LAYER VIA4 ;
    ANTENNAPARTIALCUTAREA 34.2144 LAYER T4V2 ;
    ANTENNAPARTIALCUTAREA 180.7 LAYER RV ;
    PORT
      LAYER T4M2 ;
        RECT 57 17 65 29 ;
        RECT 57 3.5 65 15.5 ;
        RECT 57 0.983 62 66.017 ;
        RECT 57 0.943 61.966 66.057 ;
        RECT 57 0.897 61.92 66.103 ;
        RECT 57 0.851 61.874 66.149 ;
        RECT 57 0.805 61.828 66.195 ;
        RECT 57 0.759 61.782 66.241 ;
        RECT 57 0.713 61.736 66.287 ;
        RECT 57 0.667 61.69 66.333 ;
        RECT 57 0.621 61.644 66.379 ;
        RECT 57 0.575 61.598 66.425 ;
        RECT 57 0.529 61.552 66.471 ;
        RECT 57 0.483 61.506 66.517 ;
        RECT 57 0.437 61.46 66.563 ;
        RECT 57 0.391 61.414 66.609 ;
        RECT 57 0.345 61.368 66.655 ;
        RECT 57 0.299 61.322 66.701 ;
        RECT 57 0.253 61.276 66.747 ;
        RECT 57 0.207 61.23 66.793 ;
        RECT 57 0.161 61.184 66.839 ;
        RECT 57 0.115 61.138 66.885 ;
        RECT 57 0.069 61.092 66.931 ;
        RECT 57 0.023 61.046 66.977 ;
        RECT 4 57.5 61 67 ;
        RECT 3 43.5 62 51 ;
        RECT 3 29.5 62 37 ;
        RECT 3 15.5 62 23 ;
        RECT 4 0 61 9 ;
        RECT 43 0 50.5 67 ;
        RECT 29 0 36.5 67 ;
        RECT 15 0 22.5 67 ;
        RECT 3 0.977 8.5 66.023 ;
        RECT 3.966 0.017 8.5 66.983 ;
        RECT 3.92 0.057 8.5 66.943 ;
        RECT 3.874 0.103 8.5 66.897 ;
        RECT 3.828 0.149 8.5 66.851 ;
        RECT 3.782 0.195 8.5 66.805 ;
        RECT 3.736 0.241 8.5 66.759 ;
        RECT 3.69 0.287 8.5 66.713 ;
        RECT 3.644 0.333 8.5 66.667 ;
        RECT 3.598 0.379 8.5 66.621 ;
        RECT 3.552 0.425 8.5 66.575 ;
        RECT 3.506 0.471 8.5 66.529 ;
        RECT 3.46 0.517 8.5 66.483 ;
        RECT 3.414 0.563 8.5 66.437 ;
        RECT 3.368 0.609 8.5 66.391 ;
        RECT 3.322 0.655 8.5 66.345 ;
        RECT 3.276 0.701 8.5 66.299 ;
        RECT 3.23 0.747 8.5 66.253 ;
        RECT 3.184 0.793 8.5 66.207 ;
        RECT 3.138 0.839 8.5 66.161 ;
        RECT 3.092 0.885 8.5 66.115 ;
        RECT 3.046 0.931 8.5 66.069 ;
        RECT 0 17 8.5 29 ;
        RECT 0 3.5 8.5 15.5 ;
      LAYER MET5 ;
        RECT 57 17 65 29 ;
        RECT 57 3.5 65 15.5 ;
        RECT 0 -14.445 65 -8.89 ;
        RECT 57 0.983 62 66.017 ;
        RECT 57 0.943 61.966 66.057 ;
        RECT 57 0.897 61.92 66.103 ;
        RECT 57 0.851 61.874 66.149 ;
        RECT 57 0.805 61.828 66.195 ;
        RECT 57 0.759 61.782 66.241 ;
        RECT 57 0.713 61.736 66.287 ;
        RECT 57 0.667 61.69 66.333 ;
        RECT 57 0.621 61.644 66.379 ;
        RECT 57 0.575 61.598 66.425 ;
        RECT 57 0.529 61.552 66.471 ;
        RECT 57 0.483 61.506 66.517 ;
        RECT 57 0.437 61.46 66.563 ;
        RECT 57 0.391 61.414 66.609 ;
        RECT 57 0.345 61.368 66.655 ;
        RECT 57 0.299 61.322 66.701 ;
        RECT 57 0.253 61.276 66.747 ;
        RECT 57 0.207 61.23 66.793 ;
        RECT 57 0.161 61.184 66.839 ;
        RECT 57 0.115 61.138 66.885 ;
        RECT 57 0.069 61.092 66.931 ;
        RECT 57 0.023 61.046 66.977 ;
        RECT 4 57.5 61 67 ;
        RECT 3 43.5 62 51 ;
        RECT 3 29.5 62 37 ;
        RECT 3 15.5 62 23 ;
        RECT 4 0 61 9 ;
        RECT 45.98 -14.445 56.98 9 ;
        RECT 43 0 50.5 67 ;
        RECT 33.32 -14.445 44.32 9 ;
        RECT 29 0 36.5 67 ;
        RECT 20.66 -14.445 31.66 9 ;
        RECT 15 0 22.5 67 ;
        RECT 8 -14.445 19 9 ;
        RECT 3 0.977 8.5 66.023 ;
        RECT 3.966 0.017 8.5 66.983 ;
        RECT 3.92 0.057 8.5 66.943 ;
        RECT 3.874 0.103 8.5 66.897 ;
        RECT 3.828 0.149 8.5 66.851 ;
        RECT 3.782 0.195 8.5 66.805 ;
        RECT 3.736 0.241 8.5 66.759 ;
        RECT 3.69 0.287 8.5 66.713 ;
        RECT 3.644 0.333 8.5 66.667 ;
        RECT 3.598 0.379 8.5 66.621 ;
        RECT 3.552 0.425 8.5 66.575 ;
        RECT 3.506 0.471 8.5 66.529 ;
        RECT 3.46 0.517 8.5 66.483 ;
        RECT 3.414 0.563 8.5 66.437 ;
        RECT 3.368 0.609 8.5 66.391 ;
        RECT 3.322 0.655 8.5 66.345 ;
        RECT 3.276 0.701 8.5 66.299 ;
        RECT 3.23 0.747 8.5 66.253 ;
        RECT 3.184 0.793 8.5 66.207 ;
        RECT 3.138 0.839 8.5 66.161 ;
        RECT 3.092 0.885 8.5 66.115 ;
        RECT 3.046 0.931 8.5 66.069 ;
        RECT 0 17 8.5 29 ;
        RECT 0 3.5 8.5 15.5 ;
        RECT 8 109 57 110 ;
      LAYER MET4 ;
        RECT 57 17 65 29 ;
        RECT 57 3.5 65 15.5 ;
        RECT 0 -14.445 65 -8.89 ;
        RECT 57 0.983 62 66.017 ;
        RECT 57 0.943 61.966 66.057 ;
        RECT 57 0.897 61.92 66.103 ;
        RECT 57 0.851 61.874 66.149 ;
        RECT 57 0.805 61.828 66.195 ;
        RECT 57 0.759 61.782 66.241 ;
        RECT 57 0.713 61.736 66.287 ;
        RECT 57 0.667 61.69 66.333 ;
        RECT 57 0.621 61.644 66.379 ;
        RECT 57 0.575 61.598 66.425 ;
        RECT 57 0.529 61.552 66.471 ;
        RECT 57 0.483 61.506 66.517 ;
        RECT 57 0.437 61.46 66.563 ;
        RECT 57 0.391 61.414 66.609 ;
        RECT 57 0.345 61.368 66.655 ;
        RECT 57 0.299 61.322 66.701 ;
        RECT 57 0.253 61.276 66.747 ;
        RECT 57 0.207 61.23 66.793 ;
        RECT 57 0.161 61.184 66.839 ;
        RECT 57 0.115 61.138 66.885 ;
        RECT 57 0.069 61.092 66.931 ;
        RECT 57 0.023 61.046 66.977 ;
        RECT 4 57.5 61 67 ;
        RECT 3 43.5 62 51 ;
        RECT 3 29.5 62 37 ;
        RECT 3 15.5 62 23 ;
        RECT 4 0 61 9 ;
        RECT 45.98 -14.445 56.98 9 ;
        RECT 43 0 50.5 67 ;
        RECT 33.32 -14.445 44.32 9 ;
        RECT 29 0 36.5 67 ;
        RECT 20.66 -14.445 31.66 9 ;
        RECT 15 0 22.5 67 ;
        RECT 8 -14.445 19 9 ;
        RECT 3 0.977 8.5 66.023 ;
        RECT 3.966 0.017 8.5 66.983 ;
        RECT 3.92 0.057 8.5 66.943 ;
        RECT 3.874 0.103 8.5 66.897 ;
        RECT 3.828 0.149 8.5 66.851 ;
        RECT 3.782 0.195 8.5 66.805 ;
        RECT 3.736 0.241 8.5 66.759 ;
        RECT 3.69 0.287 8.5 66.713 ;
        RECT 3.644 0.333 8.5 66.667 ;
        RECT 3.598 0.379 8.5 66.621 ;
        RECT 3.552 0.425 8.5 66.575 ;
        RECT 3.506 0.471 8.5 66.529 ;
        RECT 3.46 0.517 8.5 66.483 ;
        RECT 3.414 0.563 8.5 66.437 ;
        RECT 3.368 0.609 8.5 66.391 ;
        RECT 3.322 0.655 8.5 66.345 ;
        RECT 3.276 0.701 8.5 66.299 ;
        RECT 3.23 0.747 8.5 66.253 ;
        RECT 3.184 0.793 8.5 66.207 ;
        RECT 3.138 0.839 8.5 66.161 ;
        RECT 3.092 0.885 8.5 66.115 ;
        RECT 3.046 0.931 8.5 66.069 ;
        RECT 0 17 8.5 29 ;
        RECT 0 3.5 8.5 15.5 ;
        RECT 8 109 57 110 ;
      LAYER MET3 ;
        RECT 57 17 65 29 ;
        RECT 57 3.5 65 15.5 ;
        RECT 0 -14.445 65 -8.89 ;
        RECT 57 0.983 62 66.017 ;
        RECT 57 0.943 61.966 66.057 ;
        RECT 57 0.897 61.92 66.103 ;
        RECT 57 0.851 61.874 66.149 ;
        RECT 57 0.805 61.828 66.195 ;
        RECT 57 0.759 61.782 66.241 ;
        RECT 57 0.713 61.736 66.287 ;
        RECT 57 0.667 61.69 66.333 ;
        RECT 57 0.621 61.644 66.379 ;
        RECT 57 0.575 61.598 66.425 ;
        RECT 57 0.529 61.552 66.471 ;
        RECT 57 0.483 61.506 66.517 ;
        RECT 57 0.437 61.46 66.563 ;
        RECT 57 0.391 61.414 66.609 ;
        RECT 57 0.345 61.368 66.655 ;
        RECT 57 0.299 61.322 66.701 ;
        RECT 57 0.253 61.276 66.747 ;
        RECT 57 0.207 61.23 66.793 ;
        RECT 57 0.161 61.184 66.839 ;
        RECT 57 0.115 61.138 66.885 ;
        RECT 57 0.069 61.092 66.931 ;
        RECT 57 0.023 61.046 66.977 ;
        RECT 4 57.5 61 67 ;
        RECT 3 43.5 62 51 ;
        RECT 3 29.5 62 37 ;
        RECT 3 15.5 62 23 ;
        RECT 4 0 61 9 ;
        RECT 45.98 -14.445 56.98 9 ;
        RECT 43 0 50.5 67 ;
        RECT 33.32 -14.445 44.32 9 ;
        RECT 29 0 36.5 67 ;
        RECT 20.66 -14.445 31.66 9 ;
        RECT 15 0 22.5 67 ;
        RECT 8 -14.445 19 9 ;
        RECT 3 0.977 8.5 66.023 ;
        RECT 3.966 0.017 8.5 66.983 ;
        RECT 3.92 0.057 8.5 66.943 ;
        RECT 3.874 0.103 8.5 66.897 ;
        RECT 3.828 0.149 8.5 66.851 ;
        RECT 3.782 0.195 8.5 66.805 ;
        RECT 3.736 0.241 8.5 66.759 ;
        RECT 3.69 0.287 8.5 66.713 ;
        RECT 3.644 0.333 8.5 66.667 ;
        RECT 3.598 0.379 8.5 66.621 ;
        RECT 3.552 0.425 8.5 66.575 ;
        RECT 3.506 0.471 8.5 66.529 ;
        RECT 3.46 0.517 8.5 66.483 ;
        RECT 3.414 0.563 8.5 66.437 ;
        RECT 3.368 0.609 8.5 66.391 ;
        RECT 3.322 0.655 8.5 66.345 ;
        RECT 3.276 0.701 8.5 66.299 ;
        RECT 3.23 0.747 8.5 66.253 ;
        RECT 3.184 0.793 8.5 66.207 ;
        RECT 3.138 0.839 8.5 66.161 ;
        RECT 3.092 0.885 8.5 66.115 ;
        RECT 3.046 0.931 8.5 66.069 ;
        RECT 0 17 8.5 29 ;
        RECT 0 3.5 8.5 15.5 ;
        RECT 8 109 57 110 ;
      LAYER MET2 ;
        RECT 0 17 65 29 ;
        RECT 0 3.5 65 15.5 ;
        RECT 59.805 3.5 60.995 29 ;
        RECT 54.225 3.5 55.415 29 ;
        RECT 48.645 3.5 49.835 29 ;
        RECT 43.065 3.5 44.255 29 ;
        RECT 37.485 3.5 38.675 29 ;
        RECT 31.905 3.5 33.095 29 ;
        RECT 26.325 3.5 27.515 29 ;
        RECT 20.745 3.5 21.935 29 ;
        RECT 15.165 3.5 16.355 29 ;
        RECT 9.585 3.5 10.775 29 ;
        RECT 4.005 3.5 5.195 29 ;
        RECT 0 78.5 65 89.5 ;
        RECT 3 65 62 67 ;
        RECT 8 109 57 110 ;
        RECT 45.98 65 57 110 ;
        RECT 8 65 57 69.28 ;
        RECT 33.32 65 44.32 110 ;
        RECT 20.66 65 31.66 110 ;
        RECT 8 65 19 110 ;
    END
  END VSSIO
  OBS
    LAYER MET1 SPACING 0.09 ;
      RECT 0 -20 65 110 ;
    LAYER MET2 SPACING 0.1 ;
      RECT 57.175 67.175 65 78.325 ;
      RECT 62.175 63.675 65 78.325 ;
      RECT 0 77.175 7.825 78.325 ;
      RECT 6.675 67.175 7.825 78.325 ;
      RECT 6.175 77.152 7.825 78.325 ;
      RECT 6.635 76.695 7.825 78.325 ;
      RECT 6.221 77.106 7.825 78.325 ;
      RECT 6.589 76.738 7.825 78.325 ;
      RECT 6.267 77.06 7.825 78.325 ;
      RECT 6.543 76.784 7.825 78.325 ;
      RECT 6.313 77.014 7.825 78.325 ;
      RECT 6.497 76.83 7.825 78.325 ;
      RECT 6.359 76.968 7.825 78.325 ;
      RECT 6.451 76.876 7.825 78.325 ;
      RECT 6.405 76.922 7.825 78.325 ;
      RECT 6.635 67.175 7.825 68.805 ;
      RECT 6.589 67.175 7.825 68.762 ;
      RECT 6.543 67.175 7.825 68.716 ;
      RECT 6.497 67.175 7.825 68.67 ;
      RECT 6.451 67.175 7.825 68.624 ;
      RECT 6.405 67.175 7.825 68.578 ;
      RECT 6.359 67.175 7.825 68.532 ;
      RECT 6.313 67.175 7.825 68.486 ;
      RECT 6.267 67.175 7.825 68.44 ;
      RECT 6.221 67.175 7.825 68.394 ;
      RECT 6.175 67.175 7.825 68.348 ;
      RECT 0 67.175 7.825 68.325 ;
      RECT 0 63.675 2.825 68.325 ;
      RECT 0 63.675 65 64.825 ;
      RECT 0 107.675 7.825 110 ;
      RECT 6.675 89.675 7.825 110 ;
      RECT 6.175 107.652 7.825 110 ;
      RECT 6.635 107.195 7.825 110 ;
      RECT 6.221 107.606 7.825 110 ;
      RECT 6.589 107.238 7.825 110 ;
      RECT 6.267 107.56 7.825 110 ;
      RECT 6.543 107.284 7.825 110 ;
      RECT 6.313 107.514 7.825 110 ;
      RECT 6.497 107.33 7.825 110 ;
      RECT 6.359 107.468 7.825 110 ;
      RECT 6.451 107.376 7.825 110 ;
      RECT 6.405 107.422 7.825 110 ;
      RECT 6.635 97.695 7.825 99.805 ;
      RECT 6.589 97.738 7.825 99.762 ;
      RECT 6.543 97.784 7.825 99.716 ;
      RECT 6.497 97.83 7.825 99.67 ;
      RECT 6.451 97.876 7.825 99.624 ;
      RECT 6.405 97.922 7.825 99.578 ;
      RECT 6.359 97.968 7.825 99.532 ;
      RECT 6.313 98.014 7.825 99.486 ;
      RECT 6.267 98.06 7.825 99.44 ;
      RECT 6.221 98.106 7.825 99.394 ;
      RECT 6.175 98.152 7.825 99.348 ;
      RECT 0 98.175 7.825 99.325 ;
      RECT 6.635 89.675 7.825 91.305 ;
      RECT 6.589 89.675 7.825 91.262 ;
      RECT 6.543 89.675 7.825 91.216 ;
      RECT 6.497 89.675 7.825 91.17 ;
      RECT 6.451 89.675 7.825 91.124 ;
      RECT 6.405 89.675 7.825 91.078 ;
      RECT 6.359 89.675 7.825 91.032 ;
      RECT 6.313 89.675 7.825 90.986 ;
      RECT 6.267 89.675 7.825 90.94 ;
      RECT 6.221 89.675 7.825 90.894 ;
      RECT 6.175 89.675 7.825 90.848 ;
      RECT 0 89.675 7.825 90.825 ;
      RECT 0 -20 65 3.325 ;
      RECT 61.17 15.675 65 16.825 ;
      RECT 0 29.175 65 30.325 ;
      RECT 59.38 42.675 65 43.825 ;
      RECT 59.38 56.175 65 57.325 ;
      RECT 57.175 89.675 65 110 ;
      RECT 55.59 15.675 59.63 16.825 ;
      RECT 53.8 42.675 55.84 43.825 ;
      RECT 53.8 56.175 55.84 57.325 ;
      RECT 50.01 15.675 54.05 16.825 ;
      RECT 48.22 42.675 50.26 43.825 ;
      RECT 48.22 56.175 50.26 57.325 ;
      RECT 44.43 15.675 48.47 16.825 ;
      RECT 44.495 69.455 45.805 78.325 ;
      RECT 44.495 89.675 45.805 108.825 ;
      RECT 42.64 42.675 44.68 43.825 ;
      RECT 42.64 56.175 44.68 57.325 ;
      RECT 38.85 15.675 42.89 16.825 ;
      RECT 37.06 42.675 39.1 43.825 ;
      RECT 37.06 56.175 39.1 57.325 ;
      RECT 33.27 15.675 37.31 16.825 ;
      RECT 31.48 42.675 33.52 43.825 ;
      RECT 31.48 56.175 33.52 57.325 ;
      RECT 31.835 69.455 33.145 78.325 ;
      RECT 31.835 89.675 33.145 108.825 ;
      RECT 27.69 15.675 31.73 16.825 ;
      RECT 25.9 42.675 27.94 43.825 ;
      RECT 25.9 56.175 27.94 57.325 ;
      RECT 22.11 15.675 26.15 16.825 ;
      RECT 20.32 42.675 22.36 43.825 ;
      RECT 20.32 56.175 22.36 57.325 ;
      RECT 16.53 15.675 20.57 16.825 ;
      RECT 19.175 69.455 20.485 78.325 ;
      RECT 19.175 89.675 20.485 108.825 ;
      RECT 14.74 42.675 16.78 43.825 ;
      RECT 14.74 56.175 16.78 57.325 ;
      RECT 10.95 15.675 14.99 16.825 ;
      RECT 9.16 42.675 11.2 43.825 ;
      RECT 9.16 56.175 11.2 57.325 ;
      RECT 5.37 15.675 9.41 16.825 ;
      RECT 0 42.675 5.62 43.825 ;
      RECT 0 56.175 5.62 57.325 ;
      RECT 0 15.675 3.83 16.825 ;
    LAYER MET3 SPACING 0.1 ;
      RECT 62.175 -8.715 65 3.325 ;
      RECT 62.141 -8.715 65 0.808 ;
      RECT 62.095 -8.715 65 0.768 ;
      RECT 62.049 -8.715 65 0.722 ;
      RECT 62.003 -8.715 65 0.676 ;
      RECT 61.957 -8.715 65 0.63 ;
      RECT 61.911 -8.715 65 0.584 ;
      RECT 61.865 -8.715 65 0.538 ;
      RECT 61.819 -8.715 65 0.492 ;
      RECT 61.773 -8.715 65 0.446 ;
      RECT 61.727 -8.715 65 0.4 ;
      RECT 61.681 -8.715 65 0.354 ;
      RECT 61.635 -8.715 65 0.308 ;
      RECT 61.589 -8.715 65 0.262 ;
      RECT 61.543 -8.715 65 0.216 ;
      RECT 61.497 -8.715 65 0.17 ;
      RECT 61.451 -8.715 65 0.124 ;
      RECT 61.405 -8.715 65 0.078 ;
      RECT 61.359 -8.715 65 0.032 ;
      RECT 61.313 -8.715 65 -0.014 ;
      RECT 61.267 -8.715 65 -0.06 ;
      RECT 61.221 -8.715 65 -0.106 ;
      RECT 61.175 -8.715 65 -0.152 ;
      RECT 57.155 -8.715 65 -0.175 ;
      RECT 63.8 30.5 65 42.5 ;
      RECT 63.776 30.512 65 42.488 ;
      RECT 63.73 30.547 65 42.453 ;
      RECT 63.684 30.593 65 42.407 ;
      RECT 63.638 30.639 65 42.361 ;
      RECT 63.592 30.685 65 42.315 ;
      RECT 63.546 30.731 65 42.269 ;
      RECT 63.5 30.777 65 42.223 ;
      RECT 63.8 44 65 56 ;
      RECT 63.776 44.012 65 55.988 ;
      RECT 63.73 44.047 65 55.953 ;
      RECT 63.684 44.093 65 55.907 ;
      RECT 63.638 44.139 65 55.861 ;
      RECT 63.592 44.185 65 55.815 ;
      RECT 63.546 44.231 65 55.769 ;
      RECT 63.5 44.277 65 55.723 ;
      RECT 63.8 57.5 65 63.5 ;
      RECT 63.776 57.512 65 63.488 ;
      RECT 63.73 57.547 65 63.453 ;
      RECT 63.684 57.593 65 63.407 ;
      RECT 63.638 57.639 65 63.361 ;
      RECT 63.592 57.685 65 63.315 ;
      RECT 63.546 57.731 65 63.269 ;
      RECT 63.5 57.777 65 63.223 ;
      RECT 57.165 67.175 65 68.325 ;
      RECT 62.175 63.665 65 68.325 ;
      RECT 61.175 67.165 65 68.325 ;
      RECT 62.165 66.192 65 68.325 ;
      RECT 57.175 107.675 65 110 ;
      RECT 57.165 107.675 65 108.825 ;
      RECT 0 67.175 7.835 68.325 ;
      RECT 0 67.165 3.825 68.325 ;
      RECT 0 66.198 2.835 68.325 ;
      RECT 0 63.675 2.825 68.325 ;
      RECT 1.375 63.665 2.825 68.325 ;
      RECT 0 107.675 7.825 110 ;
      RECT 0 107.675 7.835 108.825 ;
      RECT 0 -8.715 2.825 3.325 ;
      RECT 0 -8.715 2.871 0.802 ;
      RECT 0 -8.715 2.917 0.756 ;
      RECT 0 -8.715 2.963 0.71 ;
      RECT 0 -8.715 3.009 0.664 ;
      RECT 0 -8.715 3.055 0.618 ;
      RECT 0 -8.715 3.101 0.572 ;
      RECT 0 -8.715 3.147 0.526 ;
      RECT 0 -8.715 3.193 0.48 ;
      RECT 0 -8.715 3.239 0.434 ;
      RECT 0 -8.715 3.285 0.388 ;
      RECT 0 -8.715 3.331 0.342 ;
      RECT 0 -8.715 3.377 0.296 ;
      RECT 0 -8.715 3.423 0.25 ;
      RECT 0 -8.715 3.469 0.204 ;
      RECT 0 -8.715 3.515 0.158 ;
      RECT 0 -8.715 3.561 0.112 ;
      RECT 0 -8.715 3.607 0.066 ;
      RECT 0 -8.715 3.653 0.02 ;
      RECT 0 -8.715 3.699 -0.026 ;
      RECT 0 -8.715 3.745 -0.072 ;
      RECT 0 -8.715 3.791 -0.118 ;
      RECT 0 -8.715 3.825 -0.158 ;
      RECT 0 -8.715 7.825 -0.175 ;
      RECT 1.375 29.175 2.825 30.335 ;
      RECT 0 29.175 2.825 30.325 ;
      RECT 1.375 42.665 2.825 43.835 ;
      RECT 0 42.675 2.825 43.825 ;
      RECT 1.375 56.165 2.825 57.335 ;
      RECT 0 56.175 2.825 57.325 ;
      RECT 0 -20 65 -14.62 ;
      RECT 62.175 15.675 65 16.825 ;
      RECT 62.175 29.175 65 30.335 ;
      RECT 62.175 42.665 65 43.835 ;
      RECT 62.175 56.165 65 57.335 ;
      RECT 57.165 77.175 65 78.335 ;
      RECT 0 78.5 65 89.5 ;
      RECT 57.165 89.665 65 90.825 ;
      RECT 57.165 98.175 65 99.325 ;
      RECT 50.675 29.165 56.825 29.325 ;
      RECT 53.79 42.665 55.85 43.325 ;
      RECT 53.79 56.165 55.85 57.325 ;
      RECT 44.485 77.175 45.815 78.335 ;
      RECT 44.485 89.665 45.815 90.825 ;
      RECT 44.485 98.175 45.815 99.325 ;
      RECT 44.485 107.675 45.815 108.825 ;
      RECT 44.495 -8.715 45.805 -0.175 ;
      RECT 36.675 29.165 42.825 29.325 ;
      RECT 42.63 42.665 42.825 43.325 ;
      RECT 42.63 56.165 42.825 57.325 ;
      RECT 37.05 42.665 39.11 43.325 ;
      RECT 37.05 56.165 39.11 57.325 ;
      RECT 31.825 77.175 33.155 78.335 ;
      RECT 31.825 89.665 33.155 90.825 ;
      RECT 31.825 98.175 33.155 99.325 ;
      RECT 31.825 107.675 33.155 108.825 ;
      RECT 31.835 -8.715 33.145 -0.175 ;
      RECT 22.675 29.165 28.825 29.325 ;
      RECT 25.89 42.665 27.95 43.325 ;
      RECT 25.89 56.165 27.95 57.325 ;
      RECT 19.165 77.175 20.495 78.335 ;
      RECT 19.165 89.665 20.495 90.825 ;
      RECT 19.165 98.175 20.495 99.325 ;
      RECT 19.165 107.675 20.495 108.825 ;
      RECT 19.175 -8.715 20.485 -0.175 ;
      RECT 8.675 29.165 14.825 29.325 ;
      RECT 9.15 42.665 11.21 43.325 ;
      RECT 9.15 56.165 11.21 57.325 ;
      RECT 0 77.175 7.835 78.335 ;
      RECT 0 89.665 7.835 90.825 ;
      RECT 0 98.175 7.835 99.325 ;
      RECT 0 15.675 2.825 16.825 ;
    LAYER MET4 SPACING 0.1 ;
      RECT 62.175 -8.715 65 3.325 ;
      RECT 62.141 -8.715 65 0.808 ;
      RECT 62.095 -8.715 65 0.768 ;
      RECT 62.049 -8.715 65 0.722 ;
      RECT 62.003 -8.715 65 0.676 ;
      RECT 61.957 -8.715 65 0.63 ;
      RECT 61.911 -8.715 65 0.584 ;
      RECT 61.865 -8.715 65 0.538 ;
      RECT 61.819 -8.715 65 0.492 ;
      RECT 61.773 -8.715 65 0.446 ;
      RECT 61.727 -8.715 65 0.4 ;
      RECT 61.681 -8.715 65 0.354 ;
      RECT 61.635 -8.715 65 0.308 ;
      RECT 61.589 -8.715 65 0.262 ;
      RECT 61.543 -8.715 65 0.216 ;
      RECT 61.497 -8.715 65 0.17 ;
      RECT 61.451 -8.715 65 0.124 ;
      RECT 61.405 -8.715 65 0.078 ;
      RECT 61.359 -8.715 65 0.032 ;
      RECT 61.313 -8.715 65 -0.014 ;
      RECT 61.267 -8.715 65 -0.06 ;
      RECT 61.221 -8.715 65 -0.106 ;
      RECT 61.175 -8.715 65 -0.152 ;
      RECT 57.155 -8.715 65 -0.175 ;
      RECT 0 67.175 65 68.325 ;
      RECT 62.175 29.175 65 68.325 ;
      RECT 61.175 67.152 65 68.325 ;
      RECT 62.141 66.192 65 68.325 ;
      RECT 0 67.158 3.825 68.325 ;
      RECT 0 67.118 3.791 68.325 ;
      RECT 61.221 67.106 65 68.325 ;
      RECT 62.095 66.232 65 68.325 ;
      RECT 0 67.072 3.745 68.325 ;
      RECT 61.267 67.06 65 68.325 ;
      RECT 62.049 66.278 65 68.325 ;
      RECT 0 67.026 3.699 68.325 ;
      RECT 61.313 67.014 65 68.325 ;
      RECT 62.003 66.324 65 68.325 ;
      RECT 0 66.98 3.653 68.325 ;
      RECT 61.359 66.968 65 68.325 ;
      RECT 61.957 66.37 65 68.325 ;
      RECT 0 66.934 3.607 68.325 ;
      RECT 61.405 66.922 65 68.325 ;
      RECT 61.911 66.416 65 68.325 ;
      RECT 0 66.888 3.561 68.325 ;
      RECT 61.451 66.876 65 68.325 ;
      RECT 61.865 66.462 65 68.325 ;
      RECT 0 66.842 3.515 68.325 ;
      RECT 61.497 66.83 65 68.325 ;
      RECT 61.819 66.508 65 68.325 ;
      RECT 0 66.796 3.469 68.325 ;
      RECT 61.543 66.784 65 68.325 ;
      RECT 61.773 66.554 65 68.325 ;
      RECT 0 66.75 3.423 68.325 ;
      RECT 61.589 66.738 65 68.325 ;
      RECT 61.727 66.6 65 68.325 ;
      RECT 0 66.704 3.377 68.325 ;
      RECT 61.635 66.692 65 68.325 ;
      RECT 61.681 66.646 65 68.325 ;
      RECT 0 66.658 3.331 68.325 ;
      RECT 0 66.612 3.285 68.325 ;
      RECT 0 66.566 3.239 68.325 ;
      RECT 0 66.52 3.193 68.325 ;
      RECT 0 66.474 3.147 68.325 ;
      RECT 0 66.428 3.101 68.325 ;
      RECT 0 66.382 3.055 68.325 ;
      RECT 0 66.336 3.009 68.325 ;
      RECT 0 66.29 2.963 68.325 ;
      RECT 0 66.244 2.917 68.325 ;
      RECT 0 66.198 2.871 68.325 ;
      RECT 0 63.675 2.825 68.325 ;
      RECT 1.675 29.175 2.825 68.325 ;
      RECT 1.375 63.652 2.825 68.325 ;
      RECT 1.651 63.387 2.825 68.325 ;
      RECT 1.421 63.606 2.825 68.325 ;
      RECT 1.605 63.422 2.825 68.325 ;
      RECT 1.467 63.56 2.825 68.325 ;
      RECT 1.559 63.468 2.825 68.325 ;
      RECT 1.513 63.514 2.825 68.325 ;
      RECT 1.651 55.887 2.825 57.613 ;
      RECT 1.605 55.922 2.825 57.578 ;
      RECT 1.559 55.968 2.825 57.532 ;
      RECT 1.513 56.014 2.825 57.486 ;
      RECT 1.467 56.06 2.825 57.44 ;
      RECT 1.421 56.106 2.825 57.394 ;
      RECT 1.375 56.152 2.825 57.348 ;
      RECT 0 56.175 2.825 57.325 ;
      RECT 1.651 42.387 2.825 44.113 ;
      RECT 1.605 42.422 2.825 44.078 ;
      RECT 1.559 42.468 2.825 44.032 ;
      RECT 1.513 42.514 2.825 43.986 ;
      RECT 1.467 42.56 2.825 43.94 ;
      RECT 1.421 42.606 2.825 43.894 ;
      RECT 1.375 42.652 2.825 43.848 ;
      RECT 0 42.675 2.825 43.825 ;
      RECT 1.651 29.175 2.825 30.613 ;
      RECT 1.605 29.175 2.825 30.578 ;
      RECT 1.559 29.175 2.825 30.532 ;
      RECT 1.513 29.175 2.825 30.486 ;
      RECT 1.467 29.175 2.825 30.44 ;
      RECT 1.421 29.175 2.825 30.394 ;
      RECT 1.375 29.175 2.825 30.348 ;
      RECT 0 29.175 2.825 30.325 ;
      RECT 57.175 107.675 65 110 ;
      RECT 0 107.675 7.825 110 ;
      RECT 0 107.675 65 108.825 ;
      RECT 0 -8.715 2.825 3.325 ;
      RECT 0 -8.715 2.871 0.802 ;
      RECT 0 -8.715 2.917 0.756 ;
      RECT 0 -8.715 2.963 0.71 ;
      RECT 0 -8.715 3.009 0.664 ;
      RECT 0 -8.715 3.055 0.618 ;
      RECT 0 -8.715 3.101 0.572 ;
      RECT 0 -8.715 3.147 0.526 ;
      RECT 0 -8.715 3.193 0.48 ;
      RECT 0 -8.715 3.239 0.434 ;
      RECT 0 -8.715 3.285 0.388 ;
      RECT 0 -8.715 3.331 0.342 ;
      RECT 0 -8.715 3.377 0.296 ;
      RECT 0 -8.715 3.423 0.25 ;
      RECT 0 -8.715 3.469 0.204 ;
      RECT 0 -8.715 3.515 0.158 ;
      RECT 0 -8.715 3.561 0.112 ;
      RECT 0 -8.715 3.607 0.066 ;
      RECT 0 -8.715 3.653 0.02 ;
      RECT 0 -8.715 3.699 -0.026 ;
      RECT 0 -8.715 3.745 -0.072 ;
      RECT 0 -8.715 3.791 -0.118 ;
      RECT 0 -8.715 3.825 -0.158 ;
      RECT 0 -8.715 7.825 -0.175 ;
      RECT 0 -20 65 -14.62 ;
      RECT 62.175 15.675 65 16.825 ;
      RECT 0 77.175 65 90.825 ;
      RECT 0 98.175 65 99.325 ;
      RECT 50.675 9.175 56.825 15.325 ;
      RECT 50.675 23.175 56.825 29.325 ;
      RECT 50.675 37.175 56.825 43.325 ;
      RECT 50.675 51.175 56.825 57.325 ;
      RECT 44.495 -8.715 45.805 -0.175 ;
      RECT 36.675 9.175 42.825 15.325 ;
      RECT 36.675 23.175 42.825 29.325 ;
      RECT 36.675 37.175 42.825 43.325 ;
      RECT 36.675 51.175 42.825 57.325 ;
      RECT 31.835 -8.715 33.145 -0.175 ;
      RECT 22.675 9.175 28.825 15.325 ;
      RECT 22.675 23.175 28.825 29.325 ;
      RECT 22.675 37.175 28.825 43.325 ;
      RECT 22.675 51.175 28.825 57.325 ;
      RECT 19.175 -8.715 20.485 -0.175 ;
      RECT 8.675 9.175 14.825 15.325 ;
      RECT 8.675 23.175 14.825 29.325 ;
      RECT 8.675 37.175 14.825 43.325 ;
      RECT 8.675 51.175 14.825 57.325 ;
      RECT 0 15.675 2.825 16.825 ;
    LAYER MET5 SPACING 0.1 ;
      RECT 62.33 -8.56 65 3.17 ;
      RECT 62.296 -8.56 65 0.653 ;
      RECT 62.25 -8.56 65 0.613 ;
      RECT 62.204 -8.56 65 0.567 ;
      RECT 62.158 -8.56 65 0.521 ;
      RECT 62.112 -8.56 65 0.475 ;
      RECT 62.066 -8.56 65 0.429 ;
      RECT 62.02 -8.56 65 0.383 ;
      RECT 61.974 -8.56 65 0.337 ;
      RECT 61.928 -8.56 65 0.291 ;
      RECT 61.882 -8.56 65 0.245 ;
      RECT 61.836 -8.56 65 0.199 ;
      RECT 61.79 -8.56 65 0.153 ;
      RECT 61.744 -8.56 65 0.107 ;
      RECT 61.698 -8.56 65 0.061 ;
      RECT 61.652 -8.56 65 0.015 ;
      RECT 61.606 -8.56 65 -0.031 ;
      RECT 61.56 -8.56 65 -0.077 ;
      RECT 61.514 -8.56 65 -0.123 ;
      RECT 61.468 -8.56 65 -0.169 ;
      RECT 61.422 -8.56 65 -0.215 ;
      RECT 61.376 -8.56 65 -0.261 ;
      RECT 61.33 -8.56 65 -0.307 ;
      RECT 57.31 -8.56 65 -0.33 ;
      RECT 0 67.33 65 68.17 ;
      RECT 62.33 29.33 65 68.17 ;
      RECT 61.33 67.307 65 68.17 ;
      RECT 62.296 66.347 65 68.17 ;
      RECT 0 67.313 3.67 68.17 ;
      RECT 0 67.273 3.636 68.17 ;
      RECT 61.376 67.261 65 68.17 ;
      RECT 62.25 66.387 65 68.17 ;
      RECT 0 67.227 3.59 68.17 ;
      RECT 61.422 67.215 65 68.17 ;
      RECT 62.204 66.433 65 68.17 ;
      RECT 0 67.181 3.544 68.17 ;
      RECT 61.468 67.169 65 68.17 ;
      RECT 62.158 66.479 65 68.17 ;
      RECT 0 67.135 3.498 68.17 ;
      RECT 61.514 67.123 65 68.17 ;
      RECT 62.112 66.525 65 68.17 ;
      RECT 0 67.089 3.452 68.17 ;
      RECT 61.56 67.077 65 68.17 ;
      RECT 62.066 66.571 65 68.17 ;
      RECT 0 67.043 3.406 68.17 ;
      RECT 61.606 67.031 65 68.17 ;
      RECT 62.02 66.617 65 68.17 ;
      RECT 0 66.997 3.36 68.17 ;
      RECT 61.652 66.985 65 68.17 ;
      RECT 61.974 66.663 65 68.17 ;
      RECT 0 66.951 3.314 68.17 ;
      RECT 61.698 66.939 65 68.17 ;
      RECT 61.928 66.709 65 68.17 ;
      RECT 0 66.905 3.268 68.17 ;
      RECT 61.744 66.893 65 68.17 ;
      RECT 61.882 66.755 65 68.17 ;
      RECT 0 66.859 3.222 68.17 ;
      RECT 61.79 66.847 65 68.17 ;
      RECT 61.836 66.801 65 68.17 ;
      RECT 0 66.813 3.176 68.17 ;
      RECT 0 66.767 3.13 68.17 ;
      RECT 0 66.721 3.084 68.17 ;
      RECT 0 66.675 3.038 68.17 ;
      RECT 0 66.629 2.992 68.17 ;
      RECT 0 66.583 2.946 68.17 ;
      RECT 0 66.537 2.9 68.17 ;
      RECT 0 66.491 2.854 68.17 ;
      RECT 0 66.445 2.808 68.17 ;
      RECT 0 66.399 2.762 68.17 ;
      RECT 0 66.353 2.716 68.17 ;
      RECT 0 63.83 2.67 68.17 ;
      RECT 1.83 29.33 2.67 68.17 ;
      RECT 1.53 63.807 2.67 68.17 ;
      RECT 1.806 63.542 2.67 68.17 ;
      RECT 1.576 63.761 2.67 68.17 ;
      RECT 1.76 63.577 2.67 68.17 ;
      RECT 1.622 63.715 2.67 68.17 ;
      RECT 1.714 63.623 2.67 68.17 ;
      RECT 1.668 63.669 2.67 68.17 ;
      RECT 1.806 56.042 2.67 57.458 ;
      RECT 1.76 56.077 2.67 57.423 ;
      RECT 1.714 56.123 2.67 57.377 ;
      RECT 1.668 56.169 2.67 57.331 ;
      RECT 1.622 56.215 2.67 57.285 ;
      RECT 1.576 56.261 2.67 57.239 ;
      RECT 1.53 56.307 2.67 57.193 ;
      RECT 0 56.33 2.67 57.17 ;
      RECT 1.806 42.542 2.67 43.958 ;
      RECT 1.76 42.577 2.67 43.923 ;
      RECT 1.714 42.623 2.67 43.877 ;
      RECT 1.668 42.669 2.67 43.831 ;
      RECT 1.622 42.715 2.67 43.785 ;
      RECT 1.576 42.761 2.67 43.739 ;
      RECT 1.53 42.807 2.67 43.693 ;
      RECT 0 42.83 2.67 43.67 ;
      RECT 1.806 29.33 2.67 30.458 ;
      RECT 1.76 29.33 2.67 30.423 ;
      RECT 1.714 29.33 2.67 30.377 ;
      RECT 1.668 29.33 2.67 30.331 ;
      RECT 1.622 29.33 2.67 30.285 ;
      RECT 1.576 29.33 2.67 30.239 ;
      RECT 1.53 29.33 2.67 30.193 ;
      RECT 0 29.33 2.67 30.17 ;
      RECT 57.33 107.83 65 110 ;
      RECT 0 107.83 7.67 110 ;
      RECT 0 107.83 65 108.67 ;
      RECT 0 -8.56 2.67 3.17 ;
      RECT 0 -8.56 2.716 0.647 ;
      RECT 0 -8.56 2.762 0.601 ;
      RECT 0 -8.56 2.808 0.555 ;
      RECT 0 -8.56 2.854 0.509 ;
      RECT 0 -8.56 2.9 0.463 ;
      RECT 0 -8.56 2.946 0.417 ;
      RECT 0 -8.56 2.992 0.371 ;
      RECT 0 -8.56 3.038 0.325 ;
      RECT 0 -8.56 3.084 0.279 ;
      RECT 0 -8.56 3.13 0.233 ;
      RECT 0 -8.56 3.176 0.187 ;
      RECT 0 -8.56 3.222 0.141 ;
      RECT 0 -8.56 3.268 0.095 ;
      RECT 0 -8.56 3.314 0.049 ;
      RECT 0 -8.56 3.36 0.003 ;
      RECT 0 -8.56 3.406 -0.043 ;
      RECT 0 -8.56 3.452 -0.089 ;
      RECT 0 -8.56 3.498 -0.135 ;
      RECT 0 -8.56 3.544 -0.181 ;
      RECT 0 -8.56 3.59 -0.227 ;
      RECT 0 -8.56 3.636 -0.273 ;
      RECT 0 -8.56 3.67 -0.313 ;
      RECT 0 -8.56 7.67 -0.33 ;
      RECT 0 -20 65 -14.775 ;
      RECT 62.33 15.83 65 16.67 ;
      RECT 0 77.33 65 90.67 ;
      RECT 0 98.33 65 99.17 ;
      RECT 50.83 9.33 56.67 15.17 ;
      RECT 50.83 23.33 56.67 29.17 ;
      RECT 50.83 37.33 56.67 43.17 ;
      RECT 50.83 51.33 56.67 57.17 ;
      RECT 44.65 -8.56 45.65 -0.33 ;
      RECT 36.83 9.33 42.67 15.17 ;
      RECT 36.83 23.33 42.67 29.17 ;
      RECT 36.83 37.33 42.67 43.17 ;
      RECT 36.83 51.33 42.67 57.17 ;
      RECT 31.99 -8.56 32.99 -0.33 ;
      RECT 22.83 9.33 28.67 15.17 ;
      RECT 22.83 23.33 28.67 29.17 ;
      RECT 22.83 37.33 28.67 43.17 ;
      RECT 22.83 51.33 28.67 57.17 ;
      RECT 19.33 -8.56 20.33 -0.33 ;
      RECT 8.83 9.33 14.67 15.17 ;
      RECT 8.83 23.33 14.67 29.17 ;
      RECT 8.83 37.33 14.67 43.17 ;
      RECT 8.83 51.33 14.67 57.17 ;
      RECT 0 15.83 2.67 16.67 ;
    LAYER T4M2 SPACING 0.4 ;
      RECT 64.584 -8.29 65 -3.193 ;
      RECT 64.538 -8.29 65 -3.239 ;
      RECT 64.492 -8.29 65 -3.285 ;
      RECT 64.446 -8.29 65 -3.331 ;
      RECT 64.4 -8.29 65 -3.377 ;
      RECT 57.58 -8.29 65 -3.4 ;
      RECT 0 -8.29 0.428 -3.205 ;
      RECT 0 -8.29 0.474 -3.251 ;
      RECT 0 -8.29 0.52 -3.297 ;
      RECT 0 -8.29 0.566 -3.343 ;
      RECT 0 -8.29 0.6 -3.383 ;
      RECT 0 -8.29 7.4 -3.4 ;
      RECT 0 -20 65 -15.045 ;
      RECT 0 -14.445 65 -8.89 ;
      RECT 0 77.6 65 90.4 ;
      RECT 57.6 108.1 65 110 ;
      RECT 44.92 -8.29 45.38 -3.4 ;
      RECT 32.26 -8.29 32.72 -3.4 ;
      RECT 19.6 -8.29 20.06 -3.4 ;
      RECT 0 108.1 7.4 110 ;
    LAYER RDL SPACING 2 ;
      RECT 0 -20 65 -5 ;
      RECT 0 72 65 110 ;
      RECT 3.5 5 61.5 63 ;
  END
END P65_1233_VSSIO3

END LIBRARY
